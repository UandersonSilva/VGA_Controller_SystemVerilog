module  font_rom ( 
        input logic font_rom_clk_in,  
        input logic [10:0] font_rom_addr_in,  
        output logic [7:0] font_rom_data_out
    ); 
  
    logic [10:0] addr_reg;

    always_ff @(posedge clk)
        addr_reg <= font_rom_addr_in;

    case(addr_reg)
        11'h000: font_rom_data_out = 8'b00000000; // 0
		11'h001: font_rom_data_out = 8'b00000000; // 1
		11'h002: font_rom_data_out = 8'b00000000; // 2
		11'h003: font_rom_data_out = 8'b00000000; // 3
		11'h004: font_rom_data_out = 8'b00000000; // 4
		11'h005: font_rom_data_out = 8'b00000000; // 5
		11'h006: font_rom_data_out = 8'b00000000; // 6
		11'h007: font_rom_data_out = 8'b00000000; // 7
		11'h008: font_rom_data_out = 8'b00000000; // 8
		11'h009: font_rom_data_out = 8'b00000000; // 9
		11'h00a: font_rom_data_out = 8'b00000000; // a
		11'h00b: font_rom_data_out = 8'b00000000; // b
		11'h00c: font_rom_data_out = 8'b00000000; // c
		11'h00d: font_rom_data_out = 8'b00000000; // d
		11'h00e: font_rom_data_out = 8'b00000000; // e
		11'h00f: font_rom_data_out = 8'b00000000; // f
		// code x01
		11'h010: font_rom_data_out = 8'b00000000; // 0
		11'h011: font_rom_data_out = 8'b00000000; // 1
		11'h012: font_rom_data_out = 8'b01111110; // 2  ******
		11'h013: font_rom_data_out = 8'b10000001; // 3 *      *
		11'h014: font_rom_data_out = 8'b10100101; // 4 * *  * *
		11'h015: font_rom_data_out = 8'b10000001; // 5 *      *
		11'h016: font_rom_data_out = 8'b10000001; // 6 *      *
		11'h017: font_rom_data_out = 8'b10111101; // 7 * **** *
		11'h018: font_rom_data_out = 8'b10011001; // 8 *  **  *
		11'h019: font_rom_data_out = 8'b10000001; // 9 *      *
		11'h01a: font_rom_data_out = 8'b10000001; // a *      *
		11'h01b: font_rom_data_out = 8'b01111110; // b  ******
		11'h01c: font_rom_data_out = 8'b00000000; // c
		11'h01d: font_rom_data_out = 8'b00000000; // d
		11'h01e: font_rom_data_out = 8'b00000000; // e
		11'h01f: font_rom_data_out = 8'b00000000; // f
		// code x02
		11'h020: font_rom_data_out = 8'b00000000; // 0
		11'h021: font_rom_data_out = 8'b00000000; // 1
		11'h022: font_rom_data_out = 8'b01111110; // 2  ******
		11'h023: font_rom_data_out = 8'b11111111; // 3 ********
		11'h024: font_rom_data_out = 8'b11011011; // 4 ** ** **
		11'h025: font_rom_data_out = 8'b11111111; // 5 ********
		11'h026: font_rom_data_out = 8'b11111111; // 6 ********
		11'h027: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h028: font_rom_data_out = 8'b11100111; // 8 ***  ***
		11'h029: font_rom_data_out = 8'b11111111; // 9 ********
		11'h02a: font_rom_data_out = 8'b11111111; // a ********
		11'h02b: font_rom_data_out = 8'b01111110; // b  ******
		11'h02c: font_rom_data_out = 8'b00000000; // c
		11'h02d: font_rom_data_out = 8'b00000000; // d
		11'h02e: font_rom_data_out = 8'b00000000; // e
		11'h02f: font_rom_data_out = 8'b00000000; // f
		// code x03
		11'h030: font_rom_data_out = 8'b00000000; // 0
		11'h031: font_rom_data_out = 8'b00000000; // 1
		11'h032: font_rom_data_out = 8'b00000000; // 2
		11'h033: font_rom_data_out = 8'b00000000; // 3
		11'h034: font_rom_data_out = 8'b01101100; // 4  ** **
		11'h035: font_rom_data_out = 8'b11111110; // 5 *******
		11'h036: font_rom_data_out = 8'b11111110; // 6 *******
		11'h037: font_rom_data_out = 8'b11111110; // 7 *******
		11'h038: font_rom_data_out = 8'b11111110; // 8 *******
		11'h039: font_rom_data_out = 8'b01111100; // 9  *****
		11'h03a: font_rom_data_out = 8'b00111000; // a   ***
		11'h03b: font_rom_data_out = 8'b00010000; // b    *
		11'h03c: font_rom_data_out = 8'b00000000; // c
		11'h03d: font_rom_data_out = 8'b00000000; // d
		11'h03e: font_rom_data_out = 8'b00000000; // e
		11'h03f: font_rom_data_out = 8'b00000000; // f
		// code x04
		11'h040: font_rom_data_out = 8'b00000000; // 0
		11'h041: font_rom_data_out = 8'b00000000; // 1
		11'h042: font_rom_data_out = 8'b00000000; // 2
		11'h043: font_rom_data_out = 8'b00000000; // 3
		11'h044: font_rom_data_out = 8'b00010000; // 4    *
		11'h045: font_rom_data_out = 8'b00111000; // 5   ***
		11'h046: font_rom_data_out = 8'b01111100; // 6  *****
		11'h047: font_rom_data_out = 8'b11111110; // 7 *******
		11'h048: font_rom_data_out = 8'b01111100; // 8  *****
		11'h049: font_rom_data_out = 8'b00111000; // 9   ***
		11'h04a: font_rom_data_out = 8'b00010000; // a    *
		11'h04b: font_rom_data_out = 8'b00000000; // b
		11'h04c: font_rom_data_out = 8'b00000000; // c
		11'h04d: font_rom_data_out = 8'b00000000; // d
		11'h04e: font_rom_data_out = 8'b00000000; // e
		11'h04f: font_rom_data_out = 8'b00000000; // f
		// code x05
		11'h050: font_rom_data_out = 8'b00000000; // 0
		11'h051: font_rom_data_out = 8'b00000000; // 1
		11'h052: font_rom_data_out = 8'b00000000; // 2
		11'h053: font_rom_data_out = 8'b00011000; // 3    **
		11'h054: font_rom_data_out = 8'b00111100; // 4   ****
		11'h055: font_rom_data_out = 8'b00111100; // 5   ****
		11'h056: font_rom_data_out = 8'b11100111; // 6 ***  ***
		11'h057: font_rom_data_out = 8'b11100111; // 7 ***  ***
		11'h058: font_rom_data_out = 8'b11100111; // 8 ***  ***
		11'h059: font_rom_data_out = 8'b00011000; // 9    **
		11'h05a: font_rom_data_out = 8'b00011000; // a    **
		11'h05b: font_rom_data_out = 8'b00111100; // b   ****
		11'h05c: font_rom_data_out = 8'b00000000; // c
		11'h05d: font_rom_data_out = 8'b00000000; // d
		11'h05e: font_rom_data_out = 8'b00000000; // e
		11'h05f: font_rom_data_out = 8'b00000000; // f
		// code x06
		11'h060: font_rom_data_out = 8'b00000000; // 0
		11'h061: font_rom_data_out = 8'b00000000; // 1
		11'h062: font_rom_data_out = 8'b00000000; // 2
		11'h063: font_rom_data_out = 8'b00011000; // 3    **
		11'h064: font_rom_data_out = 8'b00111100; // 4   ****
		11'h065: font_rom_data_out = 8'b01111110; // 5  ******
		11'h066: font_rom_data_out = 8'b11111111; // 6 ********
		11'h067: font_rom_data_out = 8'b11111111; // 7 ********
		11'h068: font_rom_data_out = 8'b01111110; // 8  ******
		11'h069: font_rom_data_out = 8'b00011000; // 9    **
		11'h06a: font_rom_data_out = 8'b00011000; // a    **
		11'h06b: font_rom_data_out = 8'b00111100; // b   ****
		11'h06c: font_rom_data_out = 8'b00000000; // c
		11'h06d: font_rom_data_out = 8'b00000000; // d
		11'h06e: font_rom_data_out = 8'b00000000; // e
		11'h06f: font_rom_data_out = 8'b00000000; // f
		// code x07
		11'h070: font_rom_data_out = 8'b00000000; // 0
		11'h071: font_rom_data_out = 8'b00000000; // 1
		11'h072: font_rom_data_out = 8'b00000000; // 2
		11'h073: font_rom_data_out = 8'b00000000; // 3
		11'h074: font_rom_data_out = 8'b00000000; // 4
		11'h075: font_rom_data_out = 8'b00000000; // 5
		11'h076: font_rom_data_out = 8'b00011000; // 6    **
		11'h077: font_rom_data_out = 8'b00111100; // 7   ****
		11'h078: font_rom_data_out = 8'b00111100; // 8   ****
		11'h079: font_rom_data_out = 8'b00011000; // 9    **
		11'h07a: font_rom_data_out = 8'b00000000; // a
		11'h07b: font_rom_data_out = 8'b00000000; // b
		11'h07c: font_rom_data_out = 8'b00000000; // c
		11'h07d: font_rom_data_out = 8'b00000000; // d
		11'h07e: font_rom_data_out = 8'b00000000; // e
		11'h07f: font_rom_data_out = 8'b00000000; // f
		// code x08
		11'h080: font_rom_data_out = 8'b11111111; // 0 ********
		11'h081: font_rom_data_out = 8'b11111111; // 1 ********
		11'h082: font_rom_data_out = 8'b11111111; // 2 ********
		11'h083: font_rom_data_out = 8'b11111111; // 3 ********
		11'h084: font_rom_data_out = 8'b11111111; // 4 ********
		11'h085: font_rom_data_out = 8'b11111111; // 5 ********
		11'h086: font_rom_data_out = 8'b11100111; // 6 ***  ***
		11'h087: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h088: font_rom_data_out = 8'b11000011; // 8 **    **
		11'h089: font_rom_data_out = 8'b11100111; // 9 ***  ***
		11'h08a: font_rom_data_out = 8'b11111111; // a ********
		11'h08b: font_rom_data_out = 8'b11111111; // b ********
		11'h08c: font_rom_data_out = 8'b11111111; // c ********
		11'h08d: font_rom_data_out = 8'b11111111; // d ********
		11'h08e: font_rom_data_out = 8'b11111111; // e ********
		11'h08f: font_rom_data_out = 8'b11111111; // f ********
		// code x09
		11'h090: font_rom_data_out = 8'b00000000; // 0
		11'h091: font_rom_data_out = 8'b00000000; // 1
		11'h092: font_rom_data_out = 8'b00000000; // 2
		11'h093: font_rom_data_out = 8'b00000000; // 3
		11'h094: font_rom_data_out = 8'b00000000; // 4
		11'h095: font_rom_data_out = 8'b00111100; // 5   ****
		11'h096: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h097: font_rom_data_out = 8'b01000010; // 7  *    *
		11'h098: font_rom_data_out = 8'b01000010; // 8  *    *
		11'h099: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h09a: font_rom_data_out = 8'b00111100; // a   ****
		11'h09b: font_rom_data_out = 8'b00000000; // b
		11'h09c: font_rom_data_out = 8'b00000000; // c
		11'h09d: font_rom_data_out = 8'b00000000; // d
		11'h09e: font_rom_data_out = 8'b00000000; // e
		11'h09f: font_rom_data_out = 8'b00000000; // f
		// code x0a
		11'h0a0: font_rom_data_out = 8'b11111111; // 0 ********
		11'h0a1: font_rom_data_out = 8'b11111111; // 1 ********
		11'h0a2: font_rom_data_out = 8'b11111111; // 2 ********
		11'h0a3: font_rom_data_out = 8'b11111111; // 3 ********
		11'h0a4: font_rom_data_out = 8'b11111111; // 4 ********
		11'h0a5: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h0a6: font_rom_data_out = 8'b10011001; // 6 *  **  *
		11'h0a7: font_rom_data_out = 8'b10111101; // 7 * **** *
		11'h0a8: font_rom_data_out = 8'b10111101; // 8 * **** *
		11'h0a9: font_rom_data_out = 8'b10011001; // 9 *  **  *
		11'h0aa: font_rom_data_out = 8'b11000011; // a **    **
		11'h0ab: font_rom_data_out = 8'b11111111; // b ********
		11'h0ac: font_rom_data_out = 8'b11111111; // c ********
		11'h0ad: font_rom_data_out = 8'b11111111; // d ********
		11'h0ae: font_rom_data_out = 8'b11111111; // e ********
		11'h0af: font_rom_data_out = 8'b11111111; // f ********
		// code x0b
		11'h0b0: font_rom_data_out = 8'b00000000; // 0
		11'h0b1: font_rom_data_out = 8'b00000000; // 1
		11'h0b2: font_rom_data_out = 8'b00011110; // 2    ****
		11'h0b3: font_rom_data_out = 8'b00001110; // 3     ***
		11'h0b4: font_rom_data_out = 8'b00011010; // 4    ** *
		11'h0b5: font_rom_data_out = 8'b00110010; // 5   **  *
		11'h0b6: font_rom_data_out = 8'b01111000; // 6  ****
		11'h0b7: font_rom_data_out = 8'b11001100; // 7 **  **
		11'h0b8: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h0b9: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h0ba: font_rom_data_out = 8'b11001100; // a **  **
		11'h0bb: font_rom_data_out = 8'b01111000; // b  ****
		11'h0bc: font_rom_data_out = 8'b00000000; // c
		11'h0bd: font_rom_data_out = 8'b00000000; // d
		11'h0be: font_rom_data_out = 8'b00000000; // e
		11'h0bf: font_rom_data_out = 8'b00000000; // f
		// code x0c
		11'h0c0: font_rom_data_out = 8'b00000000; // 0
		11'h0c1: font_rom_data_out = 8'b00000000; // 1
		11'h0c2: font_rom_data_out = 8'b00111100; // 2   ****
		11'h0c3: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h0c4: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h0c5: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h0c6: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h0c7: font_rom_data_out = 8'b00111100; // 7   ****
		11'h0c8: font_rom_data_out = 8'b00011000; // 8    **
		11'h0c9: font_rom_data_out = 8'b01111110; // 9  ******
		11'h0ca: font_rom_data_out = 8'b00011000; // a    **
		11'h0cb: font_rom_data_out = 8'b00011000; // b    **
		11'h0cc: font_rom_data_out = 8'b00000000; // c
		11'h0cd: font_rom_data_out = 8'b00000000; // d
		11'h0ce: font_rom_data_out = 8'b00000000; // e
		11'h0cf: font_rom_data_out = 8'b00000000; // f
		// code x0d
		11'h0d0: font_rom_data_out = 8'b00000000; // 0
		11'h0d1: font_rom_data_out = 8'b00000000; // 1
		11'h0d2: font_rom_data_out = 8'b00111111; // 2   ******
		11'h0d3: font_rom_data_out = 8'b00110011; // 3   **  **
		11'h0d4: font_rom_data_out = 8'b00111111; // 4   ******
		11'h0d5: font_rom_data_out = 8'b00110000; // 5   **
		11'h0d6: font_rom_data_out = 8'b00110000; // 6   **
		11'h0d7: font_rom_data_out = 8'b00110000; // 7   **
		11'h0d8: font_rom_data_out = 8'b00110000; // 8   **
		11'h0d9: font_rom_data_out = 8'b01110000; // 9  ***
		11'h0da: font_rom_data_out = 8'b11110000; // a ****
		11'h0db: font_rom_data_out = 8'b11100000; // b ***
		11'h0dc: font_rom_data_out = 8'b00000000; // c
		11'h0dd: font_rom_data_out = 8'b00000000; // d
		11'h0de: font_rom_data_out = 8'b00000000; // e
		11'h0df: font_rom_data_out = 8'b00000000; // f
		// code x0e
		11'h0e0: font_rom_data_out = 8'b00000000; // 0
		11'h0e1: font_rom_data_out = 8'b00000000; // 1
		11'h0e2: font_rom_data_out = 8'b01111111; // 2  *******
		11'h0e3: font_rom_data_out = 8'b01100011; // 3  **   **
		11'h0e4: font_rom_data_out = 8'b01111111; // 4  *******
		11'h0e5: font_rom_data_out = 8'b01100011; // 5  **   **
		11'h0e6: font_rom_data_out = 8'b01100011; // 6  **   **
		11'h0e7: font_rom_data_out = 8'b01100011; // 7  **   **
		11'h0e8: font_rom_data_out = 8'b01100011; // 8  **   **
		11'h0e9: font_rom_data_out = 8'b01100111; // 9  **  ***
		11'h0ea: font_rom_data_out = 8'b11100111; // a ***  ***
		11'h0eb: font_rom_data_out = 8'b11100110; // b ***  **
		11'h0ec: font_rom_data_out = 8'b11000000; // c **
		11'h0ed: font_rom_data_out = 8'b00000000; // d
		11'h0ee: font_rom_data_out = 8'b00000000; // e
		11'h0ef: font_rom_data_out = 8'b00000000; // f
		// code x0f
		11'h0f0: font_rom_data_out = 8'b00000000; // 0
		11'h0f1: font_rom_data_out = 8'b00000000; // 1
		11'h0f2: font_rom_data_out = 8'b00000000; // 2
		11'h0f3: font_rom_data_out = 8'b00011000; // 3    **
		11'h0f4: font_rom_data_out = 8'b00011000; // 4    **
		11'h0f5: font_rom_data_out = 8'b11011011; // 5 ** ** **
		11'h0f6: font_rom_data_out = 8'b00111100; // 6   ****
		11'h0f7: font_rom_data_out = 8'b11100111; // 7 ***  ***
		11'h0f8: font_rom_data_out = 8'b00111100; // 8   ****
		11'h0f9: font_rom_data_out = 8'b11011011; // 9 ** ** **
		11'h0fa: font_rom_data_out = 8'b00011000; // a    **
		11'h0fb: font_rom_data_out = 8'b00011000; // b    **
		11'h0fc: font_rom_data_out = 8'b00000000; // c
		11'h0fd: font_rom_data_out = 8'b00000000; // d
		11'h0fe: font_rom_data_out = 8'b00000000; // e
		11'h0ff: font_rom_data_out = 8'b00000000; // f
		// code x10
		11'h100: font_rom_data_out = 8'b00000000; // 0
		11'h101: font_rom_data_out = 8'b10000000; // 1 *
		11'h102: font_rom_data_out = 8'b11000000; // 2 **
		11'h103: font_rom_data_out = 8'b11100000; // 3 ***
		11'h104: font_rom_data_out = 8'b11110000; // 4 ****
		11'h105: font_rom_data_out = 8'b11111000; // 5 *****
		11'h106: font_rom_data_out = 8'b11111110; // 6 *******
		11'h107: font_rom_data_out = 8'b11111000; // 7 *****
		11'h108: font_rom_data_out = 8'b11110000; // 8 ****
		11'h109: font_rom_data_out = 8'b11100000; // 9 ***
		11'h10a: font_rom_data_out = 8'b11000000; // a **
		11'h10b: font_rom_data_out = 8'b10000000; // b *
		11'h10c: font_rom_data_out = 8'b00000000; // c
		11'h10d: font_rom_data_out = 8'b00000000; // d
		11'h10e: font_rom_data_out = 8'b00000000; // e
		11'h10f: font_rom_data_out = 8'b00000000; // f
		// code x11
		11'h110: font_rom_data_out = 8'b00000000; // 0
		11'h111: font_rom_data_out = 8'b00000010; // 1       *
		11'h112: font_rom_data_out = 8'b00000110; // 2      **
		11'h113: font_rom_data_out = 8'b00001110; // 3     ***
		11'h114: font_rom_data_out = 8'b00011110; // 4    ****
		11'h115: font_rom_data_out = 8'b00111110; // 5   *****
		11'h116: font_rom_data_out = 8'b11111110; // 6 *******
		11'h117: font_rom_data_out = 8'b00111110; // 7   *****
		11'h118: font_rom_data_out = 8'b00011110; // 8    ****
		11'h119: font_rom_data_out = 8'b00001110; // 9     ***
		11'h11a: font_rom_data_out = 8'b00000110; // a      **
		11'h11b: font_rom_data_out = 8'b00000010; // b       *
		11'h11c: font_rom_data_out = 8'b00000000; // c
		11'h11d: font_rom_data_out = 8'b00000000; // d
		11'h11e: font_rom_data_out = 8'b00000000; // e
		11'h11f: font_rom_data_out = 8'b00000000; // f
		// code x12
		11'h120: font_rom_data_out = 8'b00000000; // 0
		11'h121: font_rom_data_out = 8'b00000000; // 1
		11'h122: font_rom_data_out = 8'b00011000; // 2    **
		11'h123: font_rom_data_out = 8'b00111100; // 3   ****
		11'h124: font_rom_data_out = 8'b01111110; // 4  ******
		11'h125: font_rom_data_out = 8'b00011000; // 5    **
		11'h126: font_rom_data_out = 8'b00011000; // 6    **
		11'h127: font_rom_data_out = 8'b00011000; // 7    **
		11'h128: font_rom_data_out = 8'b01111110; // 8  ******
		11'h129: font_rom_data_out = 8'b00111100; // 9   ****
		11'h12a: font_rom_data_out = 8'b00011000; // a    **
		11'h12b: font_rom_data_out = 8'b00000000; // b
		11'h12c: font_rom_data_out = 8'b00000000; // c
		11'h12d: font_rom_data_out = 8'b00000000; // d
		11'h12e: font_rom_data_out = 8'b00000000; // e
		11'h12f: font_rom_data_out = 8'b00000000; // f
		// code x13
		11'h130: font_rom_data_out = 8'b00000000; // 0
		11'h131: font_rom_data_out = 8'b00000000; // 1
		11'h132: font_rom_data_out = 8'b01100110; // 2  **  **
		11'h133: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h134: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h135: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h136: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h137: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h138: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h139: font_rom_data_out = 8'b00000000; // 9
		11'h13a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h13b: font_rom_data_out = 8'b01100110; // b  **  **
		11'h13c: font_rom_data_out = 8'b00000000; // c
		11'h13d: font_rom_data_out = 8'b00000000; // d
		11'h13e: font_rom_data_out = 8'b00000000; // e
		11'h13f: font_rom_data_out = 8'b00000000; // f
		// code x14
		11'h140: font_rom_data_out = 8'b00000000; // 0
		11'h141: font_rom_data_out = 8'b00000000; // 1
		11'h142: font_rom_data_out = 8'b01111111; // 2  *******
		11'h143: font_rom_data_out = 8'b11011011; // 3 ** ** **
		11'h144: font_rom_data_out = 8'b11011011; // 4 ** ** **
		11'h145: font_rom_data_out = 8'b11011011; // 5 ** ** **
		11'h146: font_rom_data_out = 8'b01111011; // 6  **** **
		11'h147: font_rom_data_out = 8'b00011011; // 7    ** **
		11'h148: font_rom_data_out = 8'b00011011; // 8    ** **
		11'h149: font_rom_data_out = 8'b00011011; // 9    ** **
		11'h14a: font_rom_data_out = 8'b00011011; // a    ** **
		11'h14b: font_rom_data_out = 8'b00011011; // b    ** **
		11'h14c: font_rom_data_out = 8'b00000000; // c
		11'h14d: font_rom_data_out = 8'b00000000; // d
		11'h14e: font_rom_data_out = 8'b00000000; // e
		11'h14f: font_rom_data_out = 8'b00000000; // f
		// code x15
		11'h150: font_rom_data_out = 8'b00000000; // 0
		11'h151: font_rom_data_out = 8'b01111100; // 1  *****
		11'h152: font_rom_data_out = 8'b11000110; // 2 **   **
		11'h153: font_rom_data_out = 8'b01100000; // 3  **
		11'h154: font_rom_data_out = 8'b00111000; // 4   ***
		11'h155: font_rom_data_out = 8'b01101100; // 5  ** **
		11'h156: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h157: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h158: font_rom_data_out = 8'b01101100; // 8  ** **
		11'h159: font_rom_data_out = 8'b00111000; // 9   ***
		11'h15a: font_rom_data_out = 8'b00001100; // a     **
		11'h15b: font_rom_data_out = 8'b11000110; // b **   **
		11'h15c: font_rom_data_out = 8'b01111100; // c  *****
		11'h15d: font_rom_data_out = 8'b00000000; // d
		11'h15e: font_rom_data_out = 8'b00000000; // e
		11'h15f: font_rom_data_out = 8'b00000000; // f
		// code x16
		11'h160: font_rom_data_out = 8'b00000000; // 0
		11'h161: font_rom_data_out = 8'b00000000; // 1
		11'h162: font_rom_data_out = 8'b00000000; // 2
		11'h163: font_rom_data_out = 8'b00000000; // 3
		11'h164: font_rom_data_out = 8'b00000000; // 4
		11'h165: font_rom_data_out = 8'b00000000; // 5
		11'h166: font_rom_data_out = 8'b00000000; // 6
		11'h167: font_rom_data_out = 8'b00000000; // 7
		11'h168: font_rom_data_out = 8'b11111110; // 8 *******
		11'h169: font_rom_data_out = 8'b11111110; // 9 *******
		11'h16a: font_rom_data_out = 8'b11111110; // a *******
		11'h16b: font_rom_data_out = 8'b11111110; // b *******
		11'h16c: font_rom_data_out = 8'b00000000; // c
		11'h16d: font_rom_data_out = 8'b00000000; // d
		11'h16e: font_rom_data_out = 8'b00000000; // e
		11'h16f: font_rom_data_out = 8'b00000000; // f
		// code x17
		11'h170: font_rom_data_out = 8'b00000000; // 0
		11'h171: font_rom_data_out = 8'b00000000; // 1
		11'h172: font_rom_data_out = 8'b00011000; // 2    **
		11'h173: font_rom_data_out = 8'b00111100; // 3   ****
		11'h174: font_rom_data_out = 8'b01111110; // 4  ******
		11'h175: font_rom_data_out = 8'b00011000; // 5    **
		11'h176: font_rom_data_out = 8'b00011000; // 6    **
		11'h177: font_rom_data_out = 8'b00011000; // 7    **
		11'h178: font_rom_data_out = 8'b01111110; // 8  ******
		11'h179: font_rom_data_out = 8'b00111100; // 9   ****
		11'h17a: font_rom_data_out = 8'b00011000; // a    **
		11'h17b: font_rom_data_out = 8'b01111110; // b  ******
		11'h17c: font_rom_data_out = 8'b00110000; // c
		11'h17d: font_rom_data_out = 8'b00000000; // d
		11'h17e: font_rom_data_out = 8'b00000000; // e
		11'h17f: font_rom_data_out = 8'b00000000; // f
		// code x18
		11'h180: font_rom_data_out = 8'b00000000; // 0
		11'h181: font_rom_data_out = 8'b00000000; // 1
		11'h182: font_rom_data_out = 8'b00011000; // 2    **
		11'h183: font_rom_data_out = 8'b00111100; // 3   ****
		11'h184: font_rom_data_out = 8'b01111110; // 4  ******
		11'h185: font_rom_data_out = 8'b00011000; // 5    **
		11'h186: font_rom_data_out = 8'b00011000; // 6    **
		11'h187: font_rom_data_out = 8'b00011000; // 7    **
		11'h188: font_rom_data_out = 8'b00011000; // 8    **
		11'h189: font_rom_data_out = 8'b00011000; // 9    **
		11'h18a: font_rom_data_out = 8'b00011000; // a    **
		11'h18b: font_rom_data_out = 8'b00011000; // b    **
		11'h18c: font_rom_data_out = 8'b00000000; // c
		11'h18d: font_rom_data_out = 8'b00000000; // d
		11'h18e: font_rom_data_out = 8'b00000000; // e
		11'h18f: font_rom_data_out = 8'b00000000; // f
		// code x19
		11'h190: font_rom_data_out = 8'b00000000; // 0
		11'h191: font_rom_data_out = 8'b00000000; // 1
		11'h192: font_rom_data_out = 8'b00011000; // 2    **
		11'h193: font_rom_data_out = 8'b00011000; // 3    **
		11'h194: font_rom_data_out = 8'b00011000; // 4    **
		11'h195: font_rom_data_out = 8'b00011000; // 5    **
		11'h196: font_rom_data_out = 8'b00011000; // 6    **
		11'h197: font_rom_data_out = 8'b00011000; // 7    **
		11'h198: font_rom_data_out = 8'b00011000; // 8    **
		11'h199: font_rom_data_out = 8'b01111110; // 9  ******
		11'h19a: font_rom_data_out = 8'b00111100; // a   ****
		11'h19b: font_rom_data_out = 8'b00011000; // b    **
		11'h19c: font_rom_data_out = 8'b00000000; // c
		11'h19d: font_rom_data_out = 8'b00000000; // d
		11'h19e: font_rom_data_out = 8'b00000000; // e
		11'h19f: font_rom_data_out = 8'b00000000; // f
		// code x1a
		11'h1a0: font_rom_data_out = 8'b00000000; // 0
		11'h1a1: font_rom_data_out = 8'b00000000; // 1
		11'h1a2: font_rom_data_out = 8'b00000000; // 2
		11'h1a3: font_rom_data_out = 8'b00000000; // 3
		11'h1a4: font_rom_data_out = 8'b00000000; // 4
		11'h1a5: font_rom_data_out = 8'b00011000; // 5    **
		11'h1a6: font_rom_data_out = 8'b00001100; // 6     **
		11'h1a7: font_rom_data_out = 8'b11111110; // 7 *******
		11'h1a8: font_rom_data_out = 8'b00001100; // 8     **
		11'h1a9: font_rom_data_out = 8'b00011000; // 9    **
		11'h1aa: font_rom_data_out = 8'b00000000; // a
		11'h1ab: font_rom_data_out = 8'b00000000; // b
		11'h1ac: font_rom_data_out = 8'b00000000; // c
		11'h1ad: font_rom_data_out = 8'b00000000; // d
		11'h1ae: font_rom_data_out = 8'b00000000; // e
		11'h1af: font_rom_data_out = 8'b00000000; // f
		// code x1b
		11'h1b0: font_rom_data_out = 8'b00000000; // 0
		11'h1b1: font_rom_data_out = 8'b00000000; // 1
		11'h1b2: font_rom_data_out = 8'b00000000; // 2
		11'h1b3: font_rom_data_out = 8'b00000000; // 3
		11'h1b4: font_rom_data_out = 8'b00000000; // 4
		11'h1b5: font_rom_data_out = 8'b00110000; // 5   **
		11'h1b6: font_rom_data_out = 8'b01100000; // 6  **
		11'h1b7: font_rom_data_out = 8'b11111110; // 7 *******
		11'h1b8: font_rom_data_out = 8'b01100000; // 8  **
		11'h1b9: font_rom_data_out = 8'b00110000; // 9   **
		11'h1ba: font_rom_data_out = 8'b00000000; // a
		11'h1bb: font_rom_data_out = 8'b00000000; // b
		11'h1bc: font_rom_data_out = 8'b00000000; // c
		11'h1bd: font_rom_data_out = 8'b00000000; // d
		11'h1be: font_rom_data_out = 8'b00000000; // e
		11'h1bf: font_rom_data_out = 8'b00000000; // f
		// code x1c
		11'h1c0: font_rom_data_out = 8'b00000000; // 0
		11'h1c1: font_rom_data_out = 8'b00000000; // 1
		11'h1c2: font_rom_data_out = 8'b00000000; // 2
		11'h1c3: font_rom_data_out = 8'b00000000; // 3
		11'h1c4: font_rom_data_out = 8'b00000000; // 4
		11'h1c5: font_rom_data_out = 8'b00000000; // 5
		11'h1c6: font_rom_data_out = 8'b11000000; // 6 **
		11'h1c7: font_rom_data_out = 8'b11000000; // 7 **
		11'h1c8: font_rom_data_out = 8'b11000000; // 8 **
		11'h1c9: font_rom_data_out = 8'b11111110; // 9 *******
		11'h1ca: font_rom_data_out = 8'b00000000; // a
		11'h1cb: font_rom_data_out = 8'b00000000; // b
		11'h1cc: font_rom_data_out = 8'b00000000; // c
		11'h1cd: font_rom_data_out = 8'b00000000; // d
		11'h1ce: font_rom_data_out = 8'b00000000; // e
		11'h1cf: font_rom_data_out = 8'b00000000; // f
		// code x1d
		11'h1d0: font_rom_data_out = 8'b00000000; // 0
		11'h1d1: font_rom_data_out = 8'b00000000; // 1
		11'h1d2: font_rom_data_out = 8'b00000000; // 2
		11'h1d3: font_rom_data_out = 8'b00000000; // 3
		11'h1d4: font_rom_data_out = 8'b00000000; // 4
		11'h1d5: font_rom_data_out = 8'b00100100; // 5   *  *
		11'h1d6: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h1d7: font_rom_data_out = 8'b11111111; // 7 ********
		11'h1d8: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h1d9: font_rom_data_out = 8'b00100100; // 9   *  *
		11'h1da: font_rom_data_out = 8'b00000000; // a
		11'h1db: font_rom_data_out = 8'b00000000; // b
		11'h1dc: font_rom_data_out = 8'b00000000; // c
		11'h1dd: font_rom_data_out = 8'b00000000; // d
		11'h1de: font_rom_data_out = 8'b00000000; // e
		11'h1df: font_rom_data_out = 8'b00000000; // f
		// code x1e
		11'h1e0: font_rom_data_out = 8'b00000000; // 0
		11'h1e1: font_rom_data_out = 8'b00000000; // 1
		11'h1e2: font_rom_data_out = 8'b00000000; // 2
		11'h1e3: font_rom_data_out = 8'b00000000; // 3
		11'h1e4: font_rom_data_out = 8'b00010000; // 4    *
		11'h1e5: font_rom_data_out = 8'b00111000; // 5   ***
		11'h1e6: font_rom_data_out = 8'b00111000; // 6   ***
		11'h1e7: font_rom_data_out = 8'b01111100; // 7  *****
		11'h1e8: font_rom_data_out = 8'b01111100; // 8  *****
		11'h1e9: font_rom_data_out = 8'b11111110; // 9 *******
		11'h1ea: font_rom_data_out = 8'b11111110; // a *******
		11'h1eb: font_rom_data_out = 8'b00000000; // b
		11'h1ec: font_rom_data_out = 8'b00000000; // c
		11'h1ed: font_rom_data_out = 8'b00000000; // d
		11'h1ee: font_rom_data_out = 8'b00000000; // e
		11'h1ef: font_rom_data_out = 8'b00000000; // f
		// code x1f
		11'h1f0: font_rom_data_out = 8'b00000000; // 0
		11'h1f1: font_rom_data_out = 8'b00000000; // 1
		11'h1f2: font_rom_data_out = 8'b00000000; // 2
		11'h1f3: font_rom_data_out = 8'b00000000; // 3
		11'h1f4: font_rom_data_out = 8'b11111110; // 4 *******
		11'h1f5: font_rom_data_out = 8'b11111110; // 5 *******
		11'h1f6: font_rom_data_out = 8'b01111100; // 6  *****
		11'h1f7: font_rom_data_out = 8'b01111100; // 7  *****
		11'h1f8: font_rom_data_out = 8'b00111000; // 8   ***
		11'h1f9: font_rom_data_out = 8'b00111000; // 9   ***
		11'h1fa: font_rom_data_out = 8'b00010000; // a    *
		11'h1fb: font_rom_data_out = 8'b00000000; // b
		11'h1fc: font_rom_data_out = 8'b00000000; // c
		11'h1fd: font_rom_data_out = 8'b00000000; // d
		11'h1fe: font_rom_data_out = 8'b00000000; // e
		11'h1ff: font_rom_data_out = 8'b00000000; // f
		// code x20
		11'h200: font_rom_data_out = 8'b00000000; // 0
		11'h201: font_rom_data_out = 8'b00000000; // 1
		11'h202: font_rom_data_out = 8'b00000000; // 2
		11'h203: font_rom_data_out = 8'b00000000; // 3
		11'h204: font_rom_data_out = 8'b00000000; // 4
		11'h205: font_rom_data_out = 8'b00000000; // 5
		11'h206: font_rom_data_out = 8'b00000000; // 6
		11'h207: font_rom_data_out = 8'b00000000; // 7
		11'h208: font_rom_data_out = 8'b00000000; // 8
		11'h209: font_rom_data_out = 8'b00000000; // 9
		11'h20a: font_rom_data_out = 8'b00000000; // a
		11'h20b: font_rom_data_out = 8'b00000000; // b
		11'h20c: font_rom_data_out = 8'b00000000; // c
		11'h20d: font_rom_data_out = 8'b00000000; // d
		11'h20e: font_rom_data_out = 8'b00000000; // e
		11'h20f: font_rom_data_out = 8'b00000000; // f
		// code x21
		11'h210: font_rom_data_out = 8'b00000000; // 0
		11'h211: font_rom_data_out = 8'b00000000; // 1
		11'h212: font_rom_data_out = 8'b00011000; // 2    **
		11'h213: font_rom_data_out = 8'b00111100; // 3   ****
		11'h214: font_rom_data_out = 8'b00111100; // 4   ****
		11'h215: font_rom_data_out = 8'b00111100; // 5   ****
		11'h216: font_rom_data_out = 8'b00011000; // 6    **
		11'h217: font_rom_data_out = 8'b00011000; // 7    **
		11'h218: font_rom_data_out = 8'b00011000; // 8    **
		11'h219: font_rom_data_out = 8'b00000000; // 9
		11'h21a: font_rom_data_out = 8'b00011000; // a    **
		11'h21b: font_rom_data_out = 8'b00011000; // b    **
		11'h21c: font_rom_data_out = 8'b00000000; // c
		11'h21d: font_rom_data_out = 8'b00000000; // d
		11'h21e: font_rom_data_out = 8'b00000000; // e
		11'h21f: font_rom_data_out = 8'b00000000; // f
		// code x22
		11'h220: font_rom_data_out = 8'b00000000; // 0
		11'h221: font_rom_data_out = 8'b01100110; // 1  **  **
		11'h222: font_rom_data_out = 8'b01100110; // 2  **  **
		11'h223: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h224: font_rom_data_out = 8'b00100100; // 4   *  *
		11'h225: font_rom_data_out = 8'b00000000; // 5
		11'h226: font_rom_data_out = 8'b00000000; // 6
		11'h227: font_rom_data_out = 8'b00000000; // 7
		11'h228: font_rom_data_out = 8'b00000000; // 8
		11'h229: font_rom_data_out = 8'b00000000; // 9
		11'h22a: font_rom_data_out = 8'b00000000; // a
		11'h22b: font_rom_data_out = 8'b00000000; // b
		11'h22c: font_rom_data_out = 8'b00000000; // c
		11'h22d: font_rom_data_out = 8'b00000000; // d
		11'h22e: font_rom_data_out = 8'b00000000; // e
		11'h22f: font_rom_data_out = 8'b00000000; // f
		// code x23
		11'h230: font_rom_data_out = 8'b00000000; // 0
		11'h231: font_rom_data_out = 8'b00000000; // 1
		11'h232: font_rom_data_out = 8'b00000000; // 2
		11'h233: font_rom_data_out = 8'b01101100; // 3  ** **
		11'h234: font_rom_data_out = 8'b01101100; // 4  ** **
		11'h235: font_rom_data_out = 8'b11111110; // 5 *******
		11'h236: font_rom_data_out = 8'b01101100; // 6  ** **
		11'h237: font_rom_data_out = 8'b01101100; // 7  ** **
		11'h238: font_rom_data_out = 8'b01101100; // 8  ** **
		11'h239: font_rom_data_out = 8'b11111110; // 9 *******
		11'h23a: font_rom_data_out = 8'b01101100; // a  ** **
		11'h23b: font_rom_data_out = 8'b01101100; // b  ** **
		11'h23c: font_rom_data_out = 8'b00000000; // c
		11'h23d: font_rom_data_out = 8'b00000000; // d
		11'h23e: font_rom_data_out = 8'b00000000; // e
		11'h23f: font_rom_data_out = 8'b00000000; // f
		// code x24
		11'h240: font_rom_data_out = 8'b00011000; // 0     **
		11'h241: font_rom_data_out = 8'b00011000; // 1     **
		11'h242: font_rom_data_out = 8'b01111100; // 2   *****
		11'h243: font_rom_data_out = 8'b11000110; // 3  **   **
		11'h244: font_rom_data_out = 8'b11000010; // 4  **    *
		11'h245: font_rom_data_out = 8'b11000000; // 5  **
		11'h246: font_rom_data_out = 8'b01111100; // 6   *****
		11'h247: font_rom_data_out = 8'b00000110; // 7       **
		11'h248: font_rom_data_out = 8'b00000110; // 8       **
		11'h249: font_rom_data_out = 8'b10000110; // 9  *    **
		11'h24a: font_rom_data_out = 8'b11000110; // a  **   **
		11'h24b: font_rom_data_out = 8'b01111100; // b   *****
		11'h24c: font_rom_data_out = 8'b00011000; // c     **
		11'h24d: font_rom_data_out = 8'b00011000; // d     **
		11'h24e: font_rom_data_out = 8'b00000000; // e
		11'h24f: font_rom_data_out = 8'b00000000; // f
		// code x25
		11'h250: font_rom_data_out = 8'b00000000; // 0
		11'h251: font_rom_data_out = 8'b00000000; // 1
		11'h252: font_rom_data_out = 8'b00000000; // 2
		11'h253: font_rom_data_out = 8'b00000000; // 3
		11'h254: font_rom_data_out = 8'b11000010; // 4 **    *
		11'h255: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h256: font_rom_data_out = 8'b00001100; // 6     **
		11'h257: font_rom_data_out = 8'b00011000; // 7    **
		11'h258: font_rom_data_out = 8'b00110000; // 8   **
		11'h259: font_rom_data_out = 8'b01100000; // 9  **
		11'h25a: font_rom_data_out = 8'b11000110; // a **   **
		11'h25b: font_rom_data_out = 8'b10000110; // b *    **
		11'h25c: font_rom_data_out = 8'b00000000; // c
		11'h25d: font_rom_data_out = 8'b00000000; // d
		11'h25e: font_rom_data_out = 8'b00000000; // e
		11'h25f: font_rom_data_out = 8'b00000000; // f
		// code x26
		11'h260: font_rom_data_out = 8'b00000000; // 0
		11'h261: font_rom_data_out = 8'b00000000; // 1
		11'h262: font_rom_data_out = 8'b00111000; // 2   ***
		11'h263: font_rom_data_out = 8'b01101100; // 3  ** **
		11'h264: font_rom_data_out = 8'b01101100; // 4  ** **
		11'h265: font_rom_data_out = 8'b00111000; // 5   ***
		11'h266: font_rom_data_out = 8'b01110110; // 6  *** **
		11'h267: font_rom_data_out = 8'b11011100; // 7 ** ***
		11'h268: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h269: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h26a: font_rom_data_out = 8'b11001100; // a **  **
		11'h26b: font_rom_data_out = 8'b01110110; // b  *** **
		11'h26c: font_rom_data_out = 8'b00000000; // c
		11'h26d: font_rom_data_out = 8'b00000000; // d
		11'h26e: font_rom_data_out = 8'b00000000; // e
		11'h26f: font_rom_data_out = 8'b00000000; // f
		// code x27
		11'h270: font_rom_data_out = 8'b00000000; // 0
		11'h271: font_rom_data_out = 8'b00110000; // 1   **
		11'h272: font_rom_data_out = 8'b00110000; // 2   **
		11'h273: font_rom_data_out = 8'b00110000; // 3   **
		11'h274: font_rom_data_out = 8'b01100000; // 4  **
		11'h275: font_rom_data_out = 8'b00000000; // 5
		11'h276: font_rom_data_out = 8'b00000000; // 6
		11'h277: font_rom_data_out = 8'b00000000; // 7
		11'h278: font_rom_data_out = 8'b00000000; // 8
		11'h279: font_rom_data_out = 8'b00000000; // 9
		11'h27a: font_rom_data_out = 8'b00000000; // a
		11'h27b: font_rom_data_out = 8'b00000000; // b
		11'h27c: font_rom_data_out = 8'b00000000; // c
		11'h27d: font_rom_data_out = 8'b00000000; // d
		11'h27e: font_rom_data_out = 8'b00000000; // e
		11'h27f: font_rom_data_out = 8'b00000000; // f
		// code x28
		11'h280: font_rom_data_out = 8'b00000000; // 0
		11'h281: font_rom_data_out = 8'b00000000; // 1
		11'h282: font_rom_data_out = 8'b00001100; // 2     **
		11'h283: font_rom_data_out = 8'b00011000; // 3    **
		11'h284: font_rom_data_out = 8'b00110000; // 4   **
		11'h285: font_rom_data_out = 8'b00110000; // 5   **
		11'h286: font_rom_data_out = 8'b00110000; // 6   **
		11'h287: font_rom_data_out = 8'b00110000; // 7   **
		11'h288: font_rom_data_out = 8'b00110000; // 8   **
		11'h289: font_rom_data_out = 8'b00110000; // 9   **
		11'h28a: font_rom_data_out = 8'b00011000; // a    **
		11'h28b: font_rom_data_out = 8'b00001100; // b     **
		11'h28c: font_rom_data_out = 8'b00000000; // c
		11'h28d: font_rom_data_out = 8'b00000000; // d
		11'h28e: font_rom_data_out = 8'b00000000; // e
		11'h28f: font_rom_data_out = 8'b00000000; // f
		// code x29
		11'h290: font_rom_data_out = 8'b00000000; // 0
		11'h291: font_rom_data_out = 8'b00000000; // 1
		11'h292: font_rom_data_out = 8'b00110000; // 2   **
		11'h293: font_rom_data_out = 8'b00011000; // 3    **
		11'h294: font_rom_data_out = 8'b00001100; // 4     **
		11'h295: font_rom_data_out = 8'b00001100; // 5     **
		11'h296: font_rom_data_out = 8'b00001100; // 6     **
		11'h297: font_rom_data_out = 8'b00001100; // 7     **
		11'h298: font_rom_data_out = 8'b00001100; // 8     **
		11'h299: font_rom_data_out = 8'b00001100; // 9     **
		11'h29a: font_rom_data_out = 8'b00011000; // a    **
		11'h29b: font_rom_data_out = 8'b00110000; // b   **
		11'h29c: font_rom_data_out = 8'b00000000; // c
		11'h29d: font_rom_data_out = 8'b00000000; // d
		11'h29e: font_rom_data_out = 8'b00000000; // e
		11'h29f: font_rom_data_out = 8'b00000000; // f
		// code x2a
		11'h2a0: font_rom_data_out = 8'b00000000; // 0
		11'h2a1: font_rom_data_out = 8'b00000000; // 1
		11'h2a2: font_rom_data_out = 8'b00000000; // 2
		11'h2a3: font_rom_data_out = 8'b00000000; // 3
		11'h2a4: font_rom_data_out = 8'b00000000; // 4
		11'h2a5: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h2a6: font_rom_data_out = 8'b00111100; // 6   ****
		11'h2a7: font_rom_data_out = 8'b11111111; // 7 ********
		11'h2a8: font_rom_data_out = 8'b00111100; // 8   ****
		11'h2a9: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h2aa: font_rom_data_out = 8'b00000000; // a
		11'h2ab: font_rom_data_out = 8'b00000000; // b
		11'h2ac: font_rom_data_out = 8'b00000000; // c
		11'h2ad: font_rom_data_out = 8'b00000000; // d
		11'h2ae: font_rom_data_out = 8'b00000000; // e
		11'h2af: font_rom_data_out = 8'b00000000; // f
		// code x2b
		11'h2b0: font_rom_data_out = 8'b00000000; // 0
		11'h2b1: font_rom_data_out = 8'b00000000; // 1
		11'h2b2: font_rom_data_out = 8'b00000000; // 2
		11'h2b3: font_rom_data_out = 8'b00000000; // 3
		11'h2b4: font_rom_data_out = 8'b00000000; // 4
		11'h2b5: font_rom_data_out = 8'b00011000; // 5    **
		11'h2b6: font_rom_data_out = 8'b00011000; // 6    **
		11'h2b7: font_rom_data_out = 8'b01111110; // 7  ******
		11'h2b8: font_rom_data_out = 8'b00011000; // 8    **
		11'h2b9: font_rom_data_out = 8'b00011000; // 9    **
		11'h2ba: font_rom_data_out = 8'b00000000; // a
		11'h2bb: font_rom_data_out = 8'b00000000; // b
		11'h2bc: font_rom_data_out = 8'b00000000; // c
		11'h2bd: font_rom_data_out = 8'b00000000; // d
		11'h2be: font_rom_data_out = 8'b00000000; // e
		11'h2bf: font_rom_data_out = 8'b00000000; // f
		// code x2c
		11'h2c0: font_rom_data_out = 8'b00000000; // 0
		11'h2c1: font_rom_data_out = 8'b00000000; // 1
		11'h2c2: font_rom_data_out = 8'b00000000; // 2
		11'h2c3: font_rom_data_out = 8'b00000000; // 3
		11'h2c4: font_rom_data_out = 8'b00000000; // 4
		11'h2c5: font_rom_data_out = 8'b00000000; // 5
		11'h2c6: font_rom_data_out = 8'b00000000; // 6
		11'h2c7: font_rom_data_out = 8'b00000000; // 7
		11'h2c8: font_rom_data_out = 8'b00000000; // 8
		11'h2c9: font_rom_data_out = 8'b00011000; // 9    **
		11'h2ca: font_rom_data_out = 8'b00011000; // a    **
		11'h2cb: font_rom_data_out = 8'b00011000; // b    **
		11'h2cc: font_rom_data_out = 8'b00110000; // c   **
		11'h2cd: font_rom_data_out = 8'b00000000; // d
		11'h2ce: font_rom_data_out = 8'b00000000; // e
		11'h2cf: font_rom_data_out = 8'b00000000; // f
		// code x2d
		11'h2d0: font_rom_data_out = 8'b00000000; // 0
		11'h2d1: font_rom_data_out = 8'b00000000; // 1
		11'h2d2: font_rom_data_out = 8'b00000000; // 2
		11'h2d3: font_rom_data_out = 8'b00000000; // 3
		11'h2d4: font_rom_data_out = 8'b00000000; // 4
		11'h2d5: font_rom_data_out = 8'b00000000; // 5
		11'h2d6: font_rom_data_out = 8'b00000000; // 6
		11'h2d7: font_rom_data_out = 8'b01111110; // 7  ******
		11'h2d8: font_rom_data_out = 8'b00000000; // 8
		11'h2d9: font_rom_data_out = 8'b00000000; // 9
		11'h2da: font_rom_data_out = 8'b00000000; // a
		11'h2db: font_rom_data_out = 8'b00000000; // b
		11'h2dc: font_rom_data_out = 8'b00000000; // c
		11'h2dd: font_rom_data_out = 8'b00000000; // d
		11'h2de: font_rom_data_out = 8'b00000000; // e
		11'h2df: font_rom_data_out = 8'b00000000; // f
		// code x2e
		11'h2e0: font_rom_data_out = 8'b00000000; // 0
		11'h2e1: font_rom_data_out = 8'b00000000; // 1
		11'h2e2: font_rom_data_out = 8'b00000000; // 2
		11'h2e3: font_rom_data_out = 8'b00000000; // 3
		11'h2e4: font_rom_data_out = 8'b00000000; // 4
		11'h2e5: font_rom_data_out = 8'b00000000; // 5
		11'h2e6: font_rom_data_out = 8'b00000000; // 6
		11'h2e7: font_rom_data_out = 8'b00000000; // 7
		11'h2e8: font_rom_data_out = 8'b00000000; // 8
		11'h2e9: font_rom_data_out = 8'b00000000; // 9
		11'h2ea: font_rom_data_out = 8'b00011000; // a    **
		11'h2eb: font_rom_data_out = 8'b00011000; // b    **
		11'h2ec: font_rom_data_out = 8'b00000000; // c
		11'h2ed: font_rom_data_out = 8'b00000000; // d
		11'h2ee: font_rom_data_out = 8'b00000000; // e
		11'h2ef: font_rom_data_out = 8'b00000000; // f
		// code x2f
		11'h2f0: font_rom_data_out = 8'b00000000; // 0
		11'h2f1: font_rom_data_out = 8'b00000000; // 1
		11'h2f2: font_rom_data_out = 8'b00000000; // 2
		11'h2f3: font_rom_data_out = 8'b00000000; // 3
		11'h2f4: font_rom_data_out = 8'b00000010; // 4       *
		11'h2f5: font_rom_data_out = 8'b00000110; // 5      **
		11'h2f6: font_rom_data_out = 8'b00001100; // 6     **
		11'h2f7: font_rom_data_out = 8'b00011000; // 7    **
		11'h2f8: font_rom_data_out = 8'b00110000; // 8   **
		11'h2f9: font_rom_data_out = 8'b01100000; // 9  **
		11'h2fa: font_rom_data_out = 8'b11000000; // a **
		11'h2fb: font_rom_data_out = 8'b10000000; // b *
		11'h2fc: font_rom_data_out = 8'b00000000; // c
		11'h2fd: font_rom_data_out = 8'b00000000; // d
		11'h2fe: font_rom_data_out = 8'b00000000; // e
		11'h2ff: font_rom_data_out = 8'b00000000; // f
		// code x30
		11'h300: font_rom_data_out = 8'b00000000; // 0
		11'h301: font_rom_data_out = 8'b00000000; // 1
		11'h302: font_rom_data_out = 8'b01111100; // 2  *****
		11'h303: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h304: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h305: font_rom_data_out = 8'b11001110; // 5 **  ***
		11'h306: font_rom_data_out = 8'b11011110; // 6 ** ****
		11'h307: font_rom_data_out = 8'b11110110; // 7 **** **
		11'h308: font_rom_data_out = 8'b11100110; // 8 ***  **
		11'h309: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h30a: font_rom_data_out = 8'b11000110; // a **   **
		11'h30b: font_rom_data_out = 8'b01111100; // b  *****
		11'h30c: font_rom_data_out = 8'b00000000; // c
		11'h30d: font_rom_data_out = 8'b00000000; // d
		11'h30e: font_rom_data_out = 8'b00000000; // e
		11'h30f: font_rom_data_out = 8'b00000000; // f
		// code x31
		11'h310: font_rom_data_out = 8'b00000000; // 0
		11'h311: font_rom_data_out = 8'b00000000; // 1
		11'h312: font_rom_data_out = 8'b00011000; // 2
		11'h313: font_rom_data_out = 8'b00111000; // 3
		11'h314: font_rom_data_out = 8'b01111000; // 4    **
		11'h315: font_rom_data_out = 8'b00011000; // 5   ***
		11'h316: font_rom_data_out = 8'b00011000; // 6  ****
		11'h317: font_rom_data_out = 8'b00011000; // 7    **
		11'h318: font_rom_data_out = 8'b00011000; // 8    **
		11'h319: font_rom_data_out = 8'b00011000; // 9    **
		11'h31a: font_rom_data_out = 8'b00011000; // a    **
		11'h31b: font_rom_data_out = 8'b01111110; // b    **
		11'h31c: font_rom_data_out = 8'b00000000; // c    **
		11'h31d: font_rom_data_out = 8'b00000000; // d  ******
		11'h31e: font_rom_data_out = 8'b00000000; // e
		11'h31f: font_rom_data_out = 8'b00000000; // f
		// code x32
		11'h320: font_rom_data_out = 8'b00000000; // 0
		11'h321: font_rom_data_out = 8'b00000000; // 1
		11'h322: font_rom_data_out = 8'b01111100; // 2  *****
		11'h323: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h324: font_rom_data_out = 8'b00000110; // 4      **
		11'h325: font_rom_data_out = 8'b00001100; // 5     **
		11'h326: font_rom_data_out = 8'b00011000; // 6    **
		11'h327: font_rom_data_out = 8'b00110000; // 7   **
		11'h328: font_rom_data_out = 8'b01100000; // 8  **
		11'h329: font_rom_data_out = 8'b11000000; // 9 **
		11'h32a: font_rom_data_out = 8'b11000110; // a **   **
		11'h32b: font_rom_data_out = 8'b11111110; // b *******
		11'h32c: font_rom_data_out = 8'b00000000; // c
		11'h32d: font_rom_data_out = 8'b00000000; // d
		11'h32e: font_rom_data_out = 8'b00000000; // e
		11'h32f: font_rom_data_out = 8'b00000000; // f
		// code x33
		11'h330: font_rom_data_out = 8'b00000000; // 0
		11'h331: font_rom_data_out = 8'b00000000; // 1
		11'h332: font_rom_data_out = 8'b01111100; // 2  *****
		11'h333: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h334: font_rom_data_out = 8'b00000110; // 4      **
		11'h335: font_rom_data_out = 8'b00000110; // 5      **
		11'h336: font_rom_data_out = 8'b00111100; // 6   ****
		11'h337: font_rom_data_out = 8'b00000110; // 7      **
		11'h338: font_rom_data_out = 8'b00000110; // 8      **
		11'h339: font_rom_data_out = 8'b00000110; // 9      **
		11'h33a: font_rom_data_out = 8'b11000110; // a **   **
		11'h33b: font_rom_data_out = 8'b01111100; // b  *****
		11'h33c: font_rom_data_out = 8'b00000000; // c
		11'h33d: font_rom_data_out = 8'b00000000; // d
		11'h33e: font_rom_data_out = 8'b00000000; // e
		11'h33f: font_rom_data_out = 8'b00000000; // f
		// code x34
		11'h340: font_rom_data_out = 8'b00000000; // 0
		11'h341: font_rom_data_out = 8'b00000000; // 1
		11'h342: font_rom_data_out = 8'b00001100; // 2     **
		11'h343: font_rom_data_out = 8'b00011100; // 3    ***
		11'h344: font_rom_data_out = 8'b00111100; // 4   ****
		11'h345: font_rom_data_out = 8'b01101100; // 5  ** **
		11'h346: font_rom_data_out = 8'b11001100; // 6 **  **
		11'h347: font_rom_data_out = 8'b11111110; // 7 *******
		11'h348: font_rom_data_out = 8'b00001100; // 8     **
		11'h349: font_rom_data_out = 8'b00001100; // 9     **
		11'h34a: font_rom_data_out = 8'b00001100; // a     **
		11'h34b: font_rom_data_out = 8'b00011110; // b    ****
		11'h34c: font_rom_data_out = 8'b00000000; // c
		11'h34d: font_rom_data_out = 8'b00000000; // d
		11'h34e: font_rom_data_out = 8'b00000000; // e
		11'h34f: font_rom_data_out = 8'b00000000; // f
		// code x35
		11'h350: font_rom_data_out = 8'b00000000; // 0
		11'h351: font_rom_data_out = 8'b00000000; // 1
		11'h352: font_rom_data_out = 8'b11111110; // 2 *******
		11'h353: font_rom_data_out = 8'b11000000; // 3 **
		11'h354: font_rom_data_out = 8'b11000000; // 4 **
		11'h355: font_rom_data_out = 8'b11000000; // 5 **
		11'h356: font_rom_data_out = 8'b11111100; // 6 ******
		11'h357: font_rom_data_out = 8'b00000110; // 7      **
		11'h358: font_rom_data_out = 8'b00000110; // 8      **
		11'h359: font_rom_data_out = 8'b00000110; // 9      **
		11'h35a: font_rom_data_out = 8'b11000110; // a **   **
		11'h35b: font_rom_data_out = 8'b01111100; // b  *****
		11'h35c: font_rom_data_out = 8'b00000000; // c
		11'h35d: font_rom_data_out = 8'b00000000; // d
		11'h35e: font_rom_data_out = 8'b00000000; // e
		11'h35f: font_rom_data_out = 8'b00000000; // f
		// code x36
		11'h360: font_rom_data_out = 8'b00000000; // 0
		11'h361: font_rom_data_out = 8'b00000000; // 1
		11'h362: font_rom_data_out = 8'b00111000; // 2   ***
		11'h363: font_rom_data_out = 8'b01100000; // 3  **
		11'h364: font_rom_data_out = 8'b11000000; // 4 **
		11'h365: font_rom_data_out = 8'b11000000; // 5 **
		11'h366: font_rom_data_out = 8'b11111100; // 6 ******
		11'h367: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h368: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h369: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h36a: font_rom_data_out = 8'b11000110; // a **   **
		11'h36b: font_rom_data_out = 8'b01111100; // b  *****
		11'h36c: font_rom_data_out = 8'b00000000; // c
		11'h36d: font_rom_data_out = 8'b00000000; // d
		11'h36e: font_rom_data_out = 8'b00000000; // e
		11'h36f: font_rom_data_out = 8'b00000000; // f
		// code x37
		11'h370: font_rom_data_out = 8'b00000000; // 0
		11'h371: font_rom_data_out = 8'b00000000; // 1
		11'h372: font_rom_data_out = 8'b11111110; // 2 *******
		11'h373: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h374: font_rom_data_out = 8'b00000110; // 4      **
		11'h375: font_rom_data_out = 8'b00000110; // 5      **
		11'h376: font_rom_data_out = 8'b00001100; // 6     **
		11'h377: font_rom_data_out = 8'b00011000; // 7    **
		11'h378: font_rom_data_out = 8'b00110000; // 8   **
		11'h379: font_rom_data_out = 8'b00110000; // 9   **
		11'h37a: font_rom_data_out = 8'b00110000; // a   **
		11'h37b: font_rom_data_out = 8'b00110000; // b   **
		11'h37c: font_rom_data_out = 8'b00000000; // c
		11'h37d: font_rom_data_out = 8'b00000000; // d
		11'h37e: font_rom_data_out = 8'b00000000; // e
		11'h37f: font_rom_data_out = 8'b00000000; // f
		// code x38
		11'h380: font_rom_data_out = 8'b00000000; // 0
		11'h381: font_rom_data_out = 8'b00000000; // 1
		11'h382: font_rom_data_out = 8'b01111100; // 2  *****
		11'h383: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h384: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h385: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h386: font_rom_data_out = 8'b01111100; // 6  *****
		11'h387: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h388: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h389: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h38a: font_rom_data_out = 8'b11000110; // a **   **
		11'h38b: font_rom_data_out = 8'b01111100; // b  *****
		11'h38c: font_rom_data_out = 8'b00000000; // c
		11'h38d: font_rom_data_out = 8'b00000000; // d
		11'h38e: font_rom_data_out = 8'b00000000; // e
		11'h38f: font_rom_data_out = 8'b00000000; // f
		// code x39
		11'h390: font_rom_data_out = 8'b00000000; // 0
		11'h391: font_rom_data_out = 8'b00000000; // 1
		11'h392: font_rom_data_out = 8'b01111100; // 2  *****
		11'h393: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h394: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h395: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h396: font_rom_data_out = 8'b01111110; // 6  ******
		11'h397: font_rom_data_out = 8'b00000110; // 7      **
		11'h398: font_rom_data_out = 8'b00000110; // 8      **
		11'h399: font_rom_data_out = 8'b00000110; // 9      **
		11'h39a: font_rom_data_out = 8'b00001100; // a     **
		11'h39b: font_rom_data_out = 8'b01111000; // b  ****
		11'h39c: font_rom_data_out = 8'b00000000; // c
		11'h39d: font_rom_data_out = 8'b00000000; // d
		11'h39e: font_rom_data_out = 8'b00000000; // e
		11'h39f: font_rom_data_out = 8'b00000000; // f
		// code x3a
		11'h3a0: font_rom_data_out = 8'b00000000; // 0
		11'h3a1: font_rom_data_out = 8'b00000000; // 1
		11'h3a2: font_rom_data_out = 8'b00000000; // 2
		11'h3a3: font_rom_data_out = 8'b00000000; // 3
		11'h3a4: font_rom_data_out = 8'b00011000; // 4    **
		11'h3a5: font_rom_data_out = 8'b00011000; // 5    **
		11'h3a6: font_rom_data_out = 8'b00000000; // 6
		11'h3a7: font_rom_data_out = 8'b00000000; // 7
		11'h3a8: font_rom_data_out = 8'b00000000; // 8
		11'h3a9: font_rom_data_out = 8'b00011000; // 9    **
		11'h3aa: font_rom_data_out = 8'b00011000; // a    **
		11'h3ab: font_rom_data_out = 8'b00000000; // b
		11'h3ac: font_rom_data_out = 8'b00000000; // c
		11'h3ad: font_rom_data_out = 8'b00000000; // d
		11'h3ae: font_rom_data_out = 8'b00000000; // e
		11'h3af: font_rom_data_out = 8'b00000000; // f
		// code x3b
		11'h3b0: font_rom_data_out = 8'b00000000; // 0
		11'h3b1: font_rom_data_out = 8'b00000000; // 1
		11'h3b2: font_rom_data_out = 8'b00000000; // 2
		11'h3b3: font_rom_data_out = 8'b00000000; // 3
		11'h3b4: font_rom_data_out = 8'b00011000; // 4    **
		11'h3b5: font_rom_data_out = 8'b00011000; // 5    **
		11'h3b6: font_rom_data_out = 8'b00000000; // 6
		11'h3b7: font_rom_data_out = 8'b00000000; // 7
		11'h3b8: font_rom_data_out = 8'b00000000; // 8
		11'h3b9: font_rom_data_out = 8'b00011000; // 9    **
		11'h3ba: font_rom_data_out = 8'b00011000; // a    **
		11'h3bb: font_rom_data_out = 8'b00110000; // b   **
		11'h3bc: font_rom_data_out = 8'b00000000; // c
		11'h3bd: font_rom_data_out = 8'b00000000; // d
		11'h3be: font_rom_data_out = 8'b00000000; // e
		11'h3bf: font_rom_data_out = 8'b00000000; // f
		// code x3c
		11'h3c0: font_rom_data_out = 8'b00000000; // 0
		11'h3c1: font_rom_data_out = 8'b00000000; // 1
		11'h3c2: font_rom_data_out = 8'b00000000; // 2
		11'h3c3: font_rom_data_out = 8'b00000110; // 3      **
		11'h3c4: font_rom_data_out = 8'b00001100; // 4     **
		11'h3c5: font_rom_data_out = 8'b00011000; // 5    **
		11'h3c6: font_rom_data_out = 8'b00110000; // 6   **
		11'h3c7: font_rom_data_out = 8'b01100000; // 7  **
		11'h3c8: font_rom_data_out = 8'b00110000; // 8   **
		11'h3c9: font_rom_data_out = 8'b00011000; // 9    **
		11'h3ca: font_rom_data_out = 8'b00001100; // a     **
		11'h3cb: font_rom_data_out = 8'b00000110; // b      **
		11'h3cc: font_rom_data_out = 8'b00000000; // c
		11'h3cd: font_rom_data_out = 8'b00000000; // d
		11'h3ce: font_rom_data_out = 8'b00000000; // e
		11'h3cf: font_rom_data_out = 8'b00000000; // f
		// code x3d
		11'h3d0: font_rom_data_out = 8'b00000000; // 0
		11'h3d1: font_rom_data_out = 8'b00000000; // 1
		11'h3d2: font_rom_data_out = 8'b00000000; // 2
		11'h3d3: font_rom_data_out = 8'b00000000; // 3
		11'h3d4: font_rom_data_out = 8'b00000000; // 4
		11'h3d5: font_rom_data_out = 8'b01111110; // 5  ******
		11'h3d6: font_rom_data_out = 8'b00000000; // 6
		11'h3d7: font_rom_data_out = 8'b00000000; // 7
		11'h3d8: font_rom_data_out = 8'b01111110; // 8  ******
		11'h3d9: font_rom_data_out = 8'b00000000; // 9
		11'h3da: font_rom_data_out = 8'b00000000; // a
		11'h3db: font_rom_data_out = 8'b00000000; // b
		11'h3dc: font_rom_data_out = 8'b00000000; // c
		11'h3dd: font_rom_data_out = 8'b00000000; // d
		11'h3de: font_rom_data_out = 8'b00000000; // e
		11'h3df: font_rom_data_out = 8'b00000000; // f
		// code x3e
		11'h3e0: font_rom_data_out = 8'b00000000; // 0
		11'h3e1: font_rom_data_out = 8'b00000000; // 1
		11'h3e2: font_rom_data_out = 8'b00000000; // 2
		11'h3e3: font_rom_data_out = 8'b01100000; // 3  **
		11'h3e4: font_rom_data_out = 8'b00110000; // 4   **
		11'h3e5: font_rom_data_out = 8'b00011000; // 5    **
		11'h3e6: font_rom_data_out = 8'b00001100; // 6     **
		11'h3e7: font_rom_data_out = 8'b00000110; // 7      **
		11'h3e8: font_rom_data_out = 8'b00001100; // 8     **
		11'h3e9: font_rom_data_out = 8'b00011000; // 9    **
		11'h3ea: font_rom_data_out = 8'b00110000; // a   **
		11'h3eb: font_rom_data_out = 8'b01100000; // b  **
		11'h3ec: font_rom_data_out = 8'b00000000; // c
		11'h3ed: font_rom_data_out = 8'b00000000; // d
		11'h3ee: font_rom_data_out = 8'b00000000; // e
		11'h3ef: font_rom_data_out = 8'b00000000; // f
		// code x3f
		11'h3f0: font_rom_data_out = 8'b00000000; // 0
		11'h3f1: font_rom_data_out = 8'b00000000; // 1
		11'h3f2: font_rom_data_out = 8'b01111100; // 2  *****
		11'h3f3: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h3f4: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h3f5: font_rom_data_out = 8'b00001100; // 5     **
		11'h3f6: font_rom_data_out = 8'b00011000; // 6    **
		11'h3f7: font_rom_data_out = 8'b00011000; // 7    **
		11'h3f8: font_rom_data_out = 8'b00011000; // 8    **
		11'h3f9: font_rom_data_out = 8'b00000000; // 9
		11'h3fa: font_rom_data_out = 8'b00011000; // a    **
		11'h3fb: font_rom_data_out = 8'b00011000; // b    **
		11'h3fc: font_rom_data_out = 8'b00000000; // c
		11'h3fd: font_rom_data_out = 8'b00000000; // d
		11'h3fe: font_rom_data_out = 8'b00000000; // e
		11'h3ff: font_rom_data_out = 8'b00000000; // f
		// code x40
		11'h400: font_rom_data_out = 8'b00000000; // 0
		11'h401: font_rom_data_out = 8'b00000000; // 1
		11'h402: font_rom_data_out = 8'b01111100; // 2  *****
		11'h403: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h404: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h405: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h406: font_rom_data_out = 8'b11011110; // 6 ** ****
		11'h407: font_rom_data_out = 8'b11011110; // 7 ** ****
		11'h408: font_rom_data_out = 8'b11011110; // 8 ** ****
		11'h409: font_rom_data_out = 8'b11011100; // 9 ** ***
		11'h40a: font_rom_data_out = 8'b11000000; // a **
		11'h40b: font_rom_data_out = 8'b01111100; // b  *****
		11'h40c: font_rom_data_out = 8'b00000000; // c
		11'h40d: font_rom_data_out = 8'b00000000; // d
		11'h40e: font_rom_data_out = 8'b00000000; // e
		11'h40f: font_rom_data_out = 8'b00000000; // f
		// code x41
		11'h410: font_rom_data_out = 8'b00000000; // 0
		11'h411: font_rom_data_out = 8'b00000000; // 1
		11'h412: font_rom_data_out = 8'b00010000; // 2    *
		11'h413: font_rom_data_out = 8'b00111000; // 3   ***
		11'h414: font_rom_data_out = 8'b01101100; // 4  ** **
		11'h415: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h416: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h417: font_rom_data_out = 8'b11111110; // 7 *******
		11'h418: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h419: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h41a: font_rom_data_out = 8'b11000110; // a **   **
		11'h41b: font_rom_data_out = 8'b11000110; // b **   **
		11'h41c: font_rom_data_out = 8'b00000000; // c
		11'h41d: font_rom_data_out = 8'b00000000; // d
		11'h41e: font_rom_data_out = 8'b00000000; // e
		11'h41f: font_rom_data_out = 8'b00000000; // f
		// code x42
		11'h420: font_rom_data_out = 8'b00000000; // 0
		11'h421: font_rom_data_out = 8'b00000000; // 1
		11'h422: font_rom_data_out = 8'b11111100; // 2 ******
		11'h423: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h424: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h425: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h426: font_rom_data_out = 8'b01111100; // 6  *****
		11'h427: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h428: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h429: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h42a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h42b: font_rom_data_out = 8'b11111100; // b ******
		11'h42c: font_rom_data_out = 8'b00000000; // c
		11'h42d: font_rom_data_out = 8'b00000000; // d
		11'h42e: font_rom_data_out = 8'b00000000; // e
		11'h42f: font_rom_data_out = 8'b00000000; // f
		// code x43
		11'h430: font_rom_data_out = 8'b00000000; // 0
		11'h431: font_rom_data_out = 8'b00000000; // 1
		11'h432: font_rom_data_out = 8'b00111100; // 2   ****
		11'h433: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h434: font_rom_data_out = 8'b11000010; // 4 **    *
		11'h435: font_rom_data_out = 8'b11000000; // 5 **
		11'h436: font_rom_data_out = 8'b11000000; // 6 **
		11'h437: font_rom_data_out = 8'b11000000; // 7 **
		11'h438: font_rom_data_out = 8'b11000000; // 8 **
		11'h439: font_rom_data_out = 8'b11000010; // 9 **    *
		11'h43a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h43b: font_rom_data_out = 8'b00111100; // b   ****
		11'h43c: font_rom_data_out = 8'b00000000; // c
		11'h43d: font_rom_data_out = 8'b00000000; // d
		11'h43e: font_rom_data_out = 8'b00000000; // e
		11'h43f: font_rom_data_out = 8'b00000000; // f
		// code x44
		11'h440: font_rom_data_out = 8'b00000000; // 0
		11'h441: font_rom_data_out = 8'b00000000; // 1
		11'h442: font_rom_data_out = 8'b11111000; // 2 *****
		11'h443: font_rom_data_out = 8'b01101100; // 3  ** **
		11'h444: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h445: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h446: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h447: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h448: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h449: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h44a: font_rom_data_out = 8'b01101100; // a  ** **
		11'h44b: font_rom_data_out = 8'b11111000; // b *****
		11'h44c: font_rom_data_out = 8'b00000000; // c
		11'h44d: font_rom_data_out = 8'b00000000; // d
		11'h44e: font_rom_data_out = 8'b00000000; // e
		11'h44f: font_rom_data_out = 8'b00000000; // f
		// code x45
		11'h450: font_rom_data_out = 8'b00000000; // 0
		11'h451: font_rom_data_out = 8'b00000000; // 1
		11'h452: font_rom_data_out = 8'b11111110; // 2 *******
		11'h453: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h454: font_rom_data_out = 8'b01100010; // 4  **   *
		11'h455: font_rom_data_out = 8'b01101000; // 5  ** *
		11'h456: font_rom_data_out = 8'b01111000; // 6  ****
		11'h457: font_rom_data_out = 8'b01101000; // 7  ** *
		11'h458: font_rom_data_out = 8'b01100000; // 8  **
		11'h459: font_rom_data_out = 8'b01100010; // 9  **   *
		11'h45a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h45b: font_rom_data_out = 8'b11111110; // b *******
		11'h45c: font_rom_data_out = 8'b00000000; // c
		11'h45d: font_rom_data_out = 8'b00000000; // d
		11'h45e: font_rom_data_out = 8'b00000000; // e
		11'h45f: font_rom_data_out = 8'b00000000; // f
		// code x46
		11'h460: font_rom_data_out = 8'b00000000; // 0
		11'h461: font_rom_data_out = 8'b00000000; // 1
		11'h462: font_rom_data_out = 8'b11111110; // 2 *******
		11'h463: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h464: font_rom_data_out = 8'b01100010; // 4  **   *
		11'h465: font_rom_data_out = 8'b01101000; // 5  ** *
		11'h466: font_rom_data_out = 8'b01111000; // 6  ****
		11'h467: font_rom_data_out = 8'b01101000; // 7  ** *
		11'h468: font_rom_data_out = 8'b01100000; // 8  **
		11'h469: font_rom_data_out = 8'b01100000; // 9  **
		11'h46a: font_rom_data_out = 8'b01100000; // a  **
		11'h46b: font_rom_data_out = 8'b11110000; // b ****
		11'h46c: font_rom_data_out = 8'b00000000; // c
		11'h46d: font_rom_data_out = 8'b00000000; // d
		11'h46e: font_rom_data_out = 8'b00000000; // e
		11'h46f: font_rom_data_out = 8'b00000000; // f
		// code x47
		11'h470: font_rom_data_out = 8'b00000000; // 0
		11'h471: font_rom_data_out = 8'b00000000; // 1
		11'h472: font_rom_data_out = 8'b00111100; // 2   ****
		11'h473: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h474: font_rom_data_out = 8'b11000010; // 4 **    *
		11'h475: font_rom_data_out = 8'b11000000; // 5 **
		11'h476: font_rom_data_out = 8'b11000000; // 6 **
		11'h477: font_rom_data_out = 8'b11011110; // 7 ** ****
		11'h478: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h479: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h47a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h47b: font_rom_data_out = 8'b00111010; // b   *** *
		11'h47c: font_rom_data_out = 8'b00000000; // c
		11'h47d: font_rom_data_out = 8'b00000000; // d
		11'h47e: font_rom_data_out = 8'b00000000; // e
		11'h47f: font_rom_data_out = 8'b00000000; // f
		// code x48
		11'h480: font_rom_data_out = 8'b00000000; // 0
		11'h481: font_rom_data_out = 8'b00000000; // 1
		11'h482: font_rom_data_out = 8'b11000110; // 2 **   **
		11'h483: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h484: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h485: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h486: font_rom_data_out = 8'b11111110; // 6 *******
		11'h487: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h488: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h489: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h48a: font_rom_data_out = 8'b11000110; // a **   **
		11'h48b: font_rom_data_out = 8'b11000110; // b **   **
		11'h48c: font_rom_data_out = 8'b00000000; // c
		11'h48d: font_rom_data_out = 8'b00000000; // d
		11'h48e: font_rom_data_out = 8'b00000000; // e
		11'h48f: font_rom_data_out = 8'b00000000; // f
		// code x49
		11'h490: font_rom_data_out = 8'b00000000; // 0
		11'h491: font_rom_data_out = 8'b00000000; // 1
		11'h492: font_rom_data_out = 8'b00111100; // 2   ****
		11'h493: font_rom_data_out = 8'b00011000; // 3    **
		11'h494: font_rom_data_out = 8'b00011000; // 4    **
		11'h495: font_rom_data_out = 8'b00011000; // 5    **
		11'h496: font_rom_data_out = 8'b00011000; // 6    **
		11'h497: font_rom_data_out = 8'b00011000; // 7    **
		11'h498: font_rom_data_out = 8'b00011000; // 8    **
		11'h499: font_rom_data_out = 8'b00011000; // 9    **
		11'h49a: font_rom_data_out = 8'b00011000; // a    **
		11'h49b: font_rom_data_out = 8'b00111100; // b   ****
		11'h49c: font_rom_data_out = 8'b00000000; // c
		11'h49d: font_rom_data_out = 8'b00000000; // d
		11'h49e: font_rom_data_out = 8'b00000000; // e
		11'h49f: font_rom_data_out = 8'b00000000; // f
		// code x4a
		11'h4a0: font_rom_data_out = 8'b00000000; // 0
		11'h4a1: font_rom_data_out = 8'b00000000; // 1
		11'h4a2: font_rom_data_out = 8'b00011110; // 2    ****
		11'h4a3: font_rom_data_out = 8'b00001100; // 3     **
		11'h4a4: font_rom_data_out = 8'b00001100; // 4     **
		11'h4a5: font_rom_data_out = 8'b00001100; // 5     **
		11'h4a6: font_rom_data_out = 8'b00001100; // 6     **
		11'h4a7: font_rom_data_out = 8'b00001100; // 7     **
		11'h4a8: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h4a9: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h4aa: font_rom_data_out = 8'b11001100; // a **  **
		11'h4ab: font_rom_data_out = 8'b01111000; // b  ****
		11'h4ac: font_rom_data_out = 8'b00000000; // c
		11'h4ad: font_rom_data_out = 8'b00000000; // d
		11'h4ae: font_rom_data_out = 8'b00000000; // e
		11'h4af: font_rom_data_out = 8'b00000000; // f
		// code x4b
		11'h4b0: font_rom_data_out = 8'b00000000; // 0
		11'h4b1: font_rom_data_out = 8'b00000000; // 1
		11'h4b2: font_rom_data_out = 8'b11100110; // 2 ***  **
		11'h4b3: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h4b4: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h4b5: font_rom_data_out = 8'b01101100; // 5  ** **
		11'h4b6: font_rom_data_out = 8'b01111000; // 6  ****
		11'h4b7: font_rom_data_out = 8'b01111000; // 7  ****
		11'h4b8: font_rom_data_out = 8'b01101100; // 8  ** **
		11'h4b9: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h4ba: font_rom_data_out = 8'b01100110; // a  **  **
		11'h4bb: font_rom_data_out = 8'b11100110; // b ***  **
		11'h4bc: font_rom_data_out = 8'b00000000; // c
		11'h4bd: font_rom_data_out = 8'b00000000; // d
		11'h4be: font_rom_data_out = 8'b00000000; // e
		11'h4bf: font_rom_data_out = 8'b00000000; // f
		// code x4c
		11'h4c0: font_rom_data_out = 8'b00000000; // 0
		11'h4c1: font_rom_data_out = 8'b00000000; // 1
		11'h4c2: font_rom_data_out = 8'b11110000; // 2 ****
		11'h4c3: font_rom_data_out = 8'b01100000; // 3  **
		11'h4c4: font_rom_data_out = 8'b01100000; // 4  **
		11'h4c5: font_rom_data_out = 8'b01100000; // 5  **
		11'h4c6: font_rom_data_out = 8'b01100000; // 6  **
		11'h4c7: font_rom_data_out = 8'b01100000; // 7  **
		11'h4c8: font_rom_data_out = 8'b01100000; // 8  **
		11'h4c9: font_rom_data_out = 8'b01100010; // 9  **   *
		11'h4ca: font_rom_data_out = 8'b01100110; // a  **  **
		11'h4cb: font_rom_data_out = 8'b11111110; // b *******
		11'h4cc: font_rom_data_out = 8'b00000000; // c
		11'h4cd: font_rom_data_out = 8'b00000000; // d
		11'h4ce: font_rom_data_out = 8'b00000000; // e
		11'h4cf: font_rom_data_out = 8'b00000000; // f
		// code x4d
		11'h4d0: font_rom_data_out = 8'b00000000; // 0
		11'h4d1: font_rom_data_out = 8'b00000000; // 1
		11'h4d2: font_rom_data_out = 8'b11000011; // 2 **    **
		11'h4d3: font_rom_data_out = 8'b11100111; // 3 ***  ***
		11'h4d4: font_rom_data_out = 8'b11111111; // 4 ********
		11'h4d5: font_rom_data_out = 8'b11111111; // 5 ********
		11'h4d6: font_rom_data_out = 8'b11011011; // 6 ** ** **
		11'h4d7: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h4d8: font_rom_data_out = 8'b11000011; // 8 **    **
		11'h4d9: font_rom_data_out = 8'b11000011; // 9 **    **
		11'h4da: font_rom_data_out = 8'b11000011; // a **    **
		11'h4db: font_rom_data_out = 8'b11000011; // b **    **
		11'h4dc: font_rom_data_out = 8'b00000000; // c
		11'h4dd: font_rom_data_out = 8'b00000000; // d
		11'h4de: font_rom_data_out = 8'b00000000; // e
		11'h4df: font_rom_data_out = 8'b00000000; // f
		// code x4e
		11'h4e0: font_rom_data_out = 8'b00000000; // 0
		11'h4e1: font_rom_data_out = 8'b00000000; // 1
		11'h4e2: font_rom_data_out = 8'b11000110; // 2 **   **
		11'h4e3: font_rom_data_out = 8'b11100110; // 3 ***  **
		11'h4e4: font_rom_data_out = 8'b11110110; // 4 **** **
		11'h4e5: font_rom_data_out = 8'b11111110; // 5 *******
		11'h4e6: font_rom_data_out = 8'b11011110; // 6 ** ****
		11'h4e7: font_rom_data_out = 8'b11001110; // 7 **  ***
		11'h4e8: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h4e9: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h4ea: font_rom_data_out = 8'b11000110; // a **   **
		11'h4eb: font_rom_data_out = 8'b11000110; // b **   **
		11'h4ec: font_rom_data_out = 8'b00000000; // c
		11'h4ed: font_rom_data_out = 8'b00000000; // d
		11'h4ee: font_rom_data_out = 8'b00000000; // e
		11'h4ef: font_rom_data_out = 8'b00000000; // f
		// code x4f
		11'h4f0: font_rom_data_out = 8'b00000000; // 0
		11'h4f1: font_rom_data_out = 8'b00000000; // 1
		11'h4f2: font_rom_data_out = 8'b01111100; // 2  *****
		11'h4f3: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h4f4: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h4f5: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h4f6: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h4f7: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h4f8: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h4f9: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h4fa: font_rom_data_out = 8'b11000110; // a **   **
		11'h4fb: font_rom_data_out = 8'b01111100; // b  *****
		11'h4fc: font_rom_data_out = 8'b00000000; // c
		11'h4fd: font_rom_data_out = 8'b00000000; // d
		11'h4fe: font_rom_data_out = 8'b00000000; // e
		11'h4ff: font_rom_data_out = 8'b00000000; // f
		// code x50
		11'h500: font_rom_data_out = 8'b00000000; // 0
		11'h501: font_rom_data_out = 8'b00000000; // 1
		11'h502: font_rom_data_out = 8'b11111100; // 2 ******
		11'h503: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h504: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h505: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h506: font_rom_data_out = 8'b01111100; // 6  *****
		11'h507: font_rom_data_out = 8'b01100000; // 7  **
		11'h508: font_rom_data_out = 8'b01100000; // 8  **
		11'h509: font_rom_data_out = 8'b01100000; // 9  **
		11'h50a: font_rom_data_out = 8'b01100000; // a  **
		11'h50b: font_rom_data_out = 8'b11110000; // b ****
		11'h50c: font_rom_data_out = 8'b00000000; // c
		11'h50d: font_rom_data_out = 8'b00000000; // d
		11'h50e: font_rom_data_out = 8'b00000000; // e
		11'h50f: font_rom_data_out = 8'b00000000; // f
		// code x510
		11'h510: font_rom_data_out = 8'b00000000; // 0
		11'h511: font_rom_data_out = 8'b00000000; // 1
		11'h512: font_rom_data_out = 8'b01111100; // 2  *****
		11'h513: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h514: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h515: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h516: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h517: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h518: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h519: font_rom_data_out = 8'b11010110; // 9 ** * **
		11'h51a: font_rom_data_out = 8'b11011110; // a ** ****
		11'h51b: font_rom_data_out = 8'b01111100; // b  *****
		11'h51c: font_rom_data_out = 8'b00001100; // c     **
		11'h51d: font_rom_data_out = 8'b00001110; // d     ***
		11'h51e: font_rom_data_out = 8'b00000000; // e
		11'h51f: font_rom_data_out = 8'b00000000; // f
		// code x52
		11'h520: font_rom_data_out = 8'b00000000; // 0
		11'h521: font_rom_data_out = 8'b00000000; // 1
		11'h522: font_rom_data_out = 8'b11111100; // 2 ******
		11'h523: font_rom_data_out = 8'b01100110; // 3  **  **
		11'h524: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h525: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h526: font_rom_data_out = 8'b01111100; // 6  *****
		11'h527: font_rom_data_out = 8'b01101100; // 7  ** **
		11'h528: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h529: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h52a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h52b: font_rom_data_out = 8'b11100110; // b ***  **
		11'h52c: font_rom_data_out = 8'b00000000; // c
		11'h52d: font_rom_data_out = 8'b00000000; // d
		11'h52e: font_rom_data_out = 8'b00000000; // e
		11'h52f: font_rom_data_out = 8'b00000000; // f
		// code x53
		11'h530: font_rom_data_out = 8'b00000000; // 0
		11'h531: font_rom_data_out = 8'b00000000; // 1
		11'h532: font_rom_data_out = 8'b01111100; // 2  *****
		11'h533: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h534: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h535: font_rom_data_out = 8'b01100000; // 5  **
		11'h536: font_rom_data_out = 8'b00111000; // 6   ***
		11'h537: font_rom_data_out = 8'b00001100; // 7     **
		11'h538: font_rom_data_out = 8'b00000110; // 8      **
		11'h539: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h53a: font_rom_data_out = 8'b11000110; // a **   **
		11'h53b: font_rom_data_out = 8'b01111100; // b  *****
		11'h53c: font_rom_data_out = 8'b00000000; // c
		11'h53d: font_rom_data_out = 8'b00000000; // d
		11'h53e: font_rom_data_out = 8'b00000000; // e
		11'h53f: font_rom_data_out = 8'b00000000; // f
		// code x54
		11'h540: font_rom_data_out = 8'b00000000; // 0
		11'h541: font_rom_data_out = 8'b00000000; // 1
		11'h542: font_rom_data_out = 8'b11111111; // 2 ********
		11'h543: font_rom_data_out = 8'b11011011; // 3 ** ** **
		11'h544: font_rom_data_out = 8'b10011001; // 4 *  **  *
		11'h545: font_rom_data_out = 8'b00011000; // 5    **
		11'h546: font_rom_data_out = 8'b00011000; // 6    **
		11'h547: font_rom_data_out = 8'b00011000; // 7    **
		11'h548: font_rom_data_out = 8'b00011000; // 8    **
		11'h549: font_rom_data_out = 8'b00011000; // 9    **
		11'h54a: font_rom_data_out = 8'b00011000; // a    **
		11'h54b: font_rom_data_out = 8'b00111100; // b   ****
		11'h54c: font_rom_data_out = 8'b00000000; // c
		11'h54d: font_rom_data_out = 8'b00000000; // d
		11'h54e: font_rom_data_out = 8'b00000000; // e
		11'h54f: font_rom_data_out = 8'b00000000; // f
		// code x55
		11'h550: font_rom_data_out = 8'b00000000; // 0
		11'h551: font_rom_data_out = 8'b00000000; // 1
		11'h552: font_rom_data_out = 8'b11000110; // 2 **   **
		11'h553: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h554: font_rom_data_out = 8'b11000110; // 4 **   **
		11'h555: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h556: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h557: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h558: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h559: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h55a: font_rom_data_out = 8'b11000110; // a **   **
		11'h55b: font_rom_data_out = 8'b01111100; // b  *****
		11'h55c: font_rom_data_out = 8'b00000000; // c
		11'h55d: font_rom_data_out = 8'b00000000; // d
		11'h55e: font_rom_data_out = 8'b00000000; // e
		11'h55f: font_rom_data_out = 8'b00000000; // f
		// code x56
		11'h560: font_rom_data_out = 8'b00000000; // 0
		11'h561: font_rom_data_out = 8'b00000000; // 1
		11'h562: font_rom_data_out = 8'b11000011; // 2 **    **
		11'h563: font_rom_data_out = 8'b11000011; // 3 **    **
		11'h564: font_rom_data_out = 8'b11000011; // 4 **    **
		11'h565: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h566: font_rom_data_out = 8'b11000011; // 6 **    **
		11'h567: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h568: font_rom_data_out = 8'b11000011; // 8 **    **
		11'h569: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h56a: font_rom_data_out = 8'b00111100; // a   ****
		11'h56b: font_rom_data_out = 8'b00011000; // b    **
		11'h56c: font_rom_data_out = 8'b00000000; // c
		11'h56d: font_rom_data_out = 8'b00000000; // d
		11'h56e: font_rom_data_out = 8'b00000000; // e
		11'h56f: font_rom_data_out = 8'b00000000; // f
		// code x57
		11'h570: font_rom_data_out = 8'b00000000; // 0
		11'h571: font_rom_data_out = 8'b00000000; // 1
		11'h572: font_rom_data_out = 8'b11000011; // 2 **    **
		11'h573: font_rom_data_out = 8'b11000011; // 3 **    **
		11'h574: font_rom_data_out = 8'b11000011; // 4 **    **
		11'h575: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h576: font_rom_data_out = 8'b11000011; // 6 **    **
		11'h577: font_rom_data_out = 8'b11011011; // 7 ** ** **
		11'h578: font_rom_data_out = 8'b11011011; // 8 ** ** **
		11'h579: font_rom_data_out = 8'b11111111; // 9 ********
		11'h57a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h57b: font_rom_data_out = 8'b01100110; // b  **  **
		11'h57c: font_rom_data_out = 8'b00000000; // c
		11'h57d: font_rom_data_out = 8'b00000000; // d
		11'h57e: font_rom_data_out = 8'b00000000; // e
		11'h57f: font_rom_data_out = 8'b00000000; // f

		// code x58
		11'h580: font_rom_data_out = 8'b00000000; // 0
		11'h581: font_rom_data_out = 8'b00000000; // 1
		11'h582: font_rom_data_out = 8'b11000011; // 2 **    **
		11'h583: font_rom_data_out = 8'b11000011; // 3 **    **
		11'h584: font_rom_data_out = 8'b01100110; // 4  **  **
		11'h585: font_rom_data_out = 8'b00111100; // 5   ****
		11'h586: font_rom_data_out = 8'b00011000; // 6    **
		11'h587: font_rom_data_out = 8'b00011000; // 7    **
		11'h588: font_rom_data_out = 8'b00111100; // 8   ****
		11'h589: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h58a: font_rom_data_out = 8'b11000011; // a **    **
		11'h58b: font_rom_data_out = 8'b11000011; // b **    **
		11'h58c: font_rom_data_out = 8'b00000000; // c
		11'h58d: font_rom_data_out = 8'b00000000; // d
		11'h58e: font_rom_data_out = 8'b00000000; // e
		11'h58f: font_rom_data_out = 8'b00000000; // f
		// code x59
		11'h590: font_rom_data_out = 8'b00000000; // 0
		11'h591: font_rom_data_out = 8'b00000000; // 1
		11'h592: font_rom_data_out = 8'b11000011; // 2 **    **
		11'h593: font_rom_data_out = 8'b11000011; // 3 **    **
		11'h594: font_rom_data_out = 8'b11000011; // 4 **    **
		11'h595: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h596: font_rom_data_out = 8'b00111100; // 6   ****
		11'h597: font_rom_data_out = 8'b00011000; // 7    **
		11'h598: font_rom_data_out = 8'b00011000; // 8    **
		11'h599: font_rom_data_out = 8'b00011000; // 9    **
		11'h59a: font_rom_data_out = 8'b00011000; // a    **
		11'h59b: font_rom_data_out = 8'b00111100; // b   ****
		11'h59c: font_rom_data_out = 8'b00000000; // c
		11'h59d: font_rom_data_out = 8'b00000000; // d
		11'h59e: font_rom_data_out = 8'b00000000; // e
		11'h59f: font_rom_data_out = 8'b00000000; // f
		// code x5a
		11'h5a0: font_rom_data_out = 8'b00000000; // 0
		11'h5a1: font_rom_data_out = 8'b00000000; // 1
		11'h5a2: font_rom_data_out = 8'b11111111; // 2 ********
		11'h5a3: font_rom_data_out = 8'b11000011; // 3 **    **
		11'h5a4: font_rom_data_out = 8'b10000110; // 4 *    **
		11'h5a5: font_rom_data_out = 8'b00001100; // 5     **
		11'h5a6: font_rom_data_out = 8'b00011000; // 6    **
		11'h5a7: font_rom_data_out = 8'b00110000; // 7   **
		11'h5a8: font_rom_data_out = 8'b01100000; // 8  **
		11'h5a9: font_rom_data_out = 8'b11000001; // 9 **     *
		11'h5aa: font_rom_data_out = 8'b11000011; // a **    **
		11'h5ab: font_rom_data_out = 8'b11111111; // b ********
		11'h5ac: font_rom_data_out = 8'b00000000; // c
		11'h5ad: font_rom_data_out = 8'b00000000; // d
		11'h5ae: font_rom_data_out = 8'b00000000; // e
		11'h5af: font_rom_data_out = 8'b00000000; // f
		// code x5b
		11'h5b0: font_rom_data_out = 8'b00000000; // 0
		11'h5b1: font_rom_data_out = 8'b00000000; // 1
		11'h5b2: font_rom_data_out = 8'b00111100; // 2   ****
		11'h5b3: font_rom_data_out = 8'b00110000; // 3   **
		11'h5b4: font_rom_data_out = 8'b00110000; // 4   **
		11'h5b5: font_rom_data_out = 8'b00110000; // 5   **
		11'h5b6: font_rom_data_out = 8'b00110000; // 6   **
		11'h5b7: font_rom_data_out = 8'b00110000; // 7   **
		11'h5b8: font_rom_data_out = 8'b00110000; // 8   **
		11'h5b9: font_rom_data_out = 8'b00110000; // 9   **
		11'h5ba: font_rom_data_out = 8'b00110000; // a   **
		11'h5bb: font_rom_data_out = 8'b00111100; // b   ****
		11'h5bc: font_rom_data_out = 8'b00000000; // c
		11'h5bd: font_rom_data_out = 8'b00000000; // d
		11'h5be: font_rom_data_out = 8'b00000000; // e
		11'h5bf: font_rom_data_out = 8'b00000000; // f
		// code x5c
		11'h5c0: font_rom_data_out = 8'b00000000; // 0
		11'h5c1: font_rom_data_out = 8'b00000000; // 1
		11'h5c2: font_rom_data_out = 8'b00000000; // 2
		11'h5c3: font_rom_data_out = 8'b10000000; // 3 *
		11'h5c4: font_rom_data_out = 8'b11000000; // 4 **
		11'h5c5: font_rom_data_out = 8'b11100000; // 5 ***
		11'h5c6: font_rom_data_out = 8'b01110000; // 6  ***
		11'h5c7: font_rom_data_out = 8'b00111000; // 7   ***
		11'h5c8: font_rom_data_out = 8'b00011100; // 8    ***
		11'h5c9: font_rom_data_out = 8'b00001110; // 9     ***
		11'h5ca: font_rom_data_out = 8'b00000110; // a      **
		11'h5cb: font_rom_data_out = 8'b00000010; // b       *
		11'h5cc: font_rom_data_out = 8'b00000000; // c
		11'h5cd: font_rom_data_out = 8'b00000000; // d
		11'h5ce: font_rom_data_out = 8'b00000000; // e
		11'h5cf: font_rom_data_out = 8'b00000000; // f
		// code x5d
		11'h5d0: font_rom_data_out = 8'b00000000; // 0
		11'h5d1: font_rom_data_out = 8'b00000000; // 1
		11'h5d2: font_rom_data_out = 8'b00111100; // 2   ****
		11'h5d3: font_rom_data_out = 8'b00001100; // 3     **
		11'h5d4: font_rom_data_out = 8'b00001100; // 4     **
		11'h5d5: font_rom_data_out = 8'b00001100; // 5     **
		11'h5d6: font_rom_data_out = 8'b00001100; // 6     **
		11'h5d7: font_rom_data_out = 8'b00001100; // 7     **
		11'h5d8: font_rom_data_out = 8'b00001100; // 8     **
		11'h5d9: font_rom_data_out = 8'b00001100; // 9     **
		11'h5da: font_rom_data_out = 8'b00001100; // a     **
		11'h5db: font_rom_data_out = 8'b00111100; // b   ****
		11'h5dc: font_rom_data_out = 8'b00000000; // c
		11'h5dd: font_rom_data_out = 8'b00000000; // d
		11'h5de: font_rom_data_out = 8'b00000000; // e
		11'h5df: font_rom_data_out = 8'b00000000; // f
		// code x5e
		11'h5e0: font_rom_data_out = 8'b00010000; // 0    *
		11'h5e1: font_rom_data_out = 8'b00111000; // 1   ***
		11'h5e2: font_rom_data_out = 8'b01101100; // 2  ** **
		11'h5e3: font_rom_data_out = 8'b11000110; // 3 **   **
		11'h5e4: font_rom_data_out = 8'b00000000; // 4
		11'h5e5: font_rom_data_out = 8'b00000000; // 5
		11'h5e6: font_rom_data_out = 8'b00000000; // 6
		11'h5e7: font_rom_data_out = 8'b00000000; // 7
		11'h5e8: font_rom_data_out = 8'b00000000; // 8
		11'h5e9: font_rom_data_out = 8'b00000000; // 9
		11'h5ea: font_rom_data_out = 8'b00000000; // a
		11'h5eb: font_rom_data_out = 8'b00000000; // b
		11'h5ec: font_rom_data_out = 8'b00000000; // c
		11'h5ed: font_rom_data_out = 8'b00000000; // d
		11'h5ee: font_rom_data_out = 8'b00000000; // e
		11'h5ef: font_rom_data_out = 8'b00000000; // f
		// code x5f
		11'h5f0: font_rom_data_out = 8'b00000000; // 0
		11'h5f1: font_rom_data_out = 8'b00000000; // 1
		11'h5f2: font_rom_data_out = 8'b00000000; // 2
		11'h5f3: font_rom_data_out = 8'b00000000; // 3
		11'h5f4: font_rom_data_out = 8'b00000000; // 4
		11'h5f5: font_rom_data_out = 8'b00000000; // 5
		11'h5f6: font_rom_data_out = 8'b00000000; // 6
		11'h5f7: font_rom_data_out = 8'b00000000; // 7
		11'h5f8: font_rom_data_out = 8'b00000000; // 8
		11'h5f9: font_rom_data_out = 8'b00000000; // 9
		11'h5fa: font_rom_data_out = 8'b00000000; // a
		11'h5fb: font_rom_data_out = 8'b00000000; // b
		11'h5fc: font_rom_data_out = 8'b00000000; // c
		11'h5fd: font_rom_data_out = 8'b11111111; // d ********
		11'h5fe: font_rom_data_out = 8'b00000000; // e
		11'h5ff: font_rom_data_out = 8'b00000000; // f
		// code x60
		11'h600: font_rom_data_out = 8'b00110000; // 0   **
		11'h601: font_rom_data_out = 8'b00110000; // 1   **
		11'h602: font_rom_data_out = 8'b00011000; // 2    **
		11'h603: font_rom_data_out = 8'b00000000; // 3
		11'h604: font_rom_data_out = 8'b00000000; // 4
		11'h605: font_rom_data_out = 8'b00000000; // 5
		11'h606: font_rom_data_out = 8'b00000000; // 6
		11'h607: font_rom_data_out = 8'b00000000; // 7
		11'h608: font_rom_data_out = 8'b00000000; // 8
		11'h609: font_rom_data_out = 8'b00000000; // 9
		11'h60a: font_rom_data_out = 8'b00000000; // a
		11'h60b: font_rom_data_out = 8'b00000000; // b
		11'h60c: font_rom_data_out = 8'b00000000; // c
		11'h60d: font_rom_data_out = 8'b00000000; // d
		11'h60e: font_rom_data_out = 8'b00000000; // e
		11'h60f: font_rom_data_out = 8'b00000000; // f
		// code x61
		11'h610: font_rom_data_out = 8'b00000000; // 0
		11'h611: font_rom_data_out = 8'b00000000; // 1
		11'h612: font_rom_data_out = 8'b00000000; // 2
		11'h613: font_rom_data_out = 8'b00000000; // 3
		11'h614: font_rom_data_out = 8'b00000000; // 4
		11'h615: font_rom_data_out = 8'b01111000; // 5  ****
		11'h616: font_rom_data_out = 8'b00001100; // 6     **
		11'h617: font_rom_data_out = 8'b01111100; // 7  *****
		11'h618: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h619: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h61a: font_rom_data_out = 8'b11001100; // a **  **
		11'h61b: font_rom_data_out = 8'b01110110; // b  *** **
		11'h61c: font_rom_data_out = 8'b00000000; // c
		11'h61d: font_rom_data_out = 8'b00000000; // d
		11'h61e: font_rom_data_out = 8'b00000000; // e
		11'h61f: font_rom_data_out = 8'b00000000; // f
		// code x62
		11'h620: font_rom_data_out = 8'b00000000; // 0
		11'h621: font_rom_data_out = 8'b00000000; // 1
		11'h622: font_rom_data_out = 8'b11100000; // 2  ***
		11'h623: font_rom_data_out = 8'b01100000; // 3   **
		11'h624: font_rom_data_out = 8'b01100000; // 4   **
		11'h625: font_rom_data_out = 8'b01111000; // 5   ****
		11'h626: font_rom_data_out = 8'b01101100; // 6   ** **
		11'h627: font_rom_data_out = 8'b01100110; // 7   **  **
		11'h628: font_rom_data_out = 8'b01100110; // 8   **  **
		11'h629: font_rom_data_out = 8'b01100110; // 9   **  **
		11'h62a: font_rom_data_out = 8'b01100110; // a   **  **
		11'h62b: font_rom_data_out = 8'b01111100; // b   *****
		11'h62c: font_rom_data_out = 8'b00000000; // c
		11'h62d: font_rom_data_out = 8'b00000000; // d
		11'h62e: font_rom_data_out = 8'b00000000; // e
		11'h62f: font_rom_data_out = 8'b00000000; // f
		// code x63
		11'h630: font_rom_data_out = 8'b00000000; // 0
		11'h631: font_rom_data_out = 8'b00000000; // 1
		11'h632: font_rom_data_out = 8'b00000000; // 2
		11'h633: font_rom_data_out = 8'b00000000; // 3
		11'h634: font_rom_data_out = 8'b00000000; // 4
		11'h635: font_rom_data_out = 8'b01111100; // 5  *****
		11'h636: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h637: font_rom_data_out = 8'b11000000; // 7 **
		11'h638: font_rom_data_out = 8'b11000000; // 8 **
		11'h639: font_rom_data_out = 8'b11000000; // 9 **
		11'h63a: font_rom_data_out = 8'b11000110; // a **   **
		11'h63b: font_rom_data_out = 8'b01111100; // b  *****
		11'h63c: font_rom_data_out = 8'b00000000; // c
		11'h63d: font_rom_data_out = 8'b00000000; // d
		11'h63e: font_rom_data_out = 8'b00000000; // e
		11'h63f: font_rom_data_out = 8'b00000000; // f
		// code x64
		11'h640: font_rom_data_out = 8'b00000000; // 0
		11'h641: font_rom_data_out = 8'b00000000; // 1
		11'h642: font_rom_data_out = 8'b00011100; // 2    ***
		11'h643: font_rom_data_out = 8'b00001100; // 3     **
		11'h644: font_rom_data_out = 8'b00001100; // 4     **
		11'h645: font_rom_data_out = 8'b00111100; // 5   ****
		11'h646: font_rom_data_out = 8'b01101100; // 6  ** **
		11'h647: font_rom_data_out = 8'b11001100; // 7 **  **
		11'h648: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h649: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h64a: font_rom_data_out = 8'b11001100; // a **  **
		11'h64b: font_rom_data_out = 8'b01110110; // b  *** **
		11'h64c: font_rom_data_out = 8'b00000000; // c
		11'h64d: font_rom_data_out = 8'b00000000; // d
		11'h64e: font_rom_data_out = 8'b00000000; // e
		11'h64f: font_rom_data_out = 8'b00000000; // f
		// code x65
		11'h650: font_rom_data_out = 8'b00000000; // 0
		11'h651: font_rom_data_out = 8'b00000000; // 1
		11'h652: font_rom_data_out = 8'b00000000; // 2
		11'h653: font_rom_data_out = 8'b00000000; // 3
		11'h654: font_rom_data_out = 8'b00000000; // 4
		11'h655: font_rom_data_out = 8'b01111100; // 5  *****
		11'h656: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h657: font_rom_data_out = 8'b11111110; // 7 *******
		11'h658: font_rom_data_out = 8'b11000000; // 8 **
		11'h659: font_rom_data_out = 8'b11000000; // 9 **
		11'h65a: font_rom_data_out = 8'b11000110; // a **   **
		11'h65b: font_rom_data_out = 8'b01111100; // b  *****
		11'h65c: font_rom_data_out = 8'b00000000; // c
		11'h65d: font_rom_data_out = 8'b00000000; // d
		11'h65e: font_rom_data_out = 8'b00000000; // e
		11'h65f: font_rom_data_out = 8'b00000000; // f
		// code x66
		11'h660: font_rom_data_out = 8'b00000000; // 0
		11'h661: font_rom_data_out = 8'b00000000; // 1
		11'h662: font_rom_data_out = 8'b00111000; // 2   ***
		11'h663: font_rom_data_out = 8'b01101100; // 3  ** **
		11'h664: font_rom_data_out = 8'b01100100; // 4  **  *
		11'h665: font_rom_data_out = 8'b01100000; // 5  **
		11'h666: font_rom_data_out = 8'b11110000; // 6 ****
		11'h667: font_rom_data_out = 8'b01100000; // 7  **
		11'h668: font_rom_data_out = 8'b01100000; // 8  **
		11'h669: font_rom_data_out = 8'b01100000; // 9  **
		11'h66a: font_rom_data_out = 8'b01100000; // a  **
		11'h66b: font_rom_data_out = 8'b11110000; // b ****
		11'h66c: font_rom_data_out = 8'b00000000; // c
		11'h66d: font_rom_data_out = 8'b00000000; // d
		11'h66e: font_rom_data_out = 8'b00000000; // e
		11'h66f: font_rom_data_out = 8'b00000000; // f
		// code x67
		11'h670: font_rom_data_out = 8'b00000000; // 0
		11'h671: font_rom_data_out = 8'b00000000; // 1
		11'h672: font_rom_data_out = 8'b00000000; // 2
		11'h673: font_rom_data_out = 8'b00000000; // 3
		11'h674: font_rom_data_out = 8'b00000000; // 4
		11'h675: font_rom_data_out = 8'b01110110; // 5  *** **
		11'h676: font_rom_data_out = 8'b11001100; // 6 **  **
		11'h677: font_rom_data_out = 8'b11001100; // 7 **  **
		11'h678: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h679: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h67a: font_rom_data_out = 8'b11001100; // a **  **
		11'h67b: font_rom_data_out = 8'b01111100; // b  *****
		11'h67c: font_rom_data_out = 8'b00001100; // c     **
		11'h67d: font_rom_data_out = 8'b11001100; // d **  **
		11'h67e: font_rom_data_out = 8'b01111000; // e  ****
		11'h67f: font_rom_data_out = 8'b00000000; // f
		// code x68
		11'h680: font_rom_data_out = 8'b00000000; // 0
		11'h681: font_rom_data_out = 8'b00000000; // 1
		11'h682: font_rom_data_out = 8'b11100000; // 2 ***
		11'h683: font_rom_data_out = 8'b01100000; // 3  **
		11'h684: font_rom_data_out = 8'b01100000; // 4  **
		11'h685: font_rom_data_out = 8'b01101100; // 5  ** **
		11'h686: font_rom_data_out = 8'b01110110; // 6  *** **
		11'h687: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h688: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h689: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h68a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h68b: font_rom_data_out = 8'b11100110; // b ***  **
		11'h68c: font_rom_data_out = 8'b00000000; // c
		11'h68d: font_rom_data_out = 8'b00000000; // d
		11'h68e: font_rom_data_out = 8'b00000000; // e
		11'h68f: font_rom_data_out = 8'b00000000; // f
		// code x69
		11'h690: font_rom_data_out = 8'b00000000; // 0
		11'h691: font_rom_data_out = 8'b00000000; // 1
		11'h692: font_rom_data_out = 8'b00011000; // 2    **
		11'h693: font_rom_data_out = 8'b00011000; // 3    **
		11'h694: font_rom_data_out = 8'b00000000; // 4
		11'h695: font_rom_data_out = 8'b00111000; // 5   ***
		11'h696: font_rom_data_out = 8'b00011000; // 6    **
		11'h697: font_rom_data_out = 8'b00011000; // 7    **
		11'h698: font_rom_data_out = 8'b00011000; // 8    **
		11'h699: font_rom_data_out = 8'b00011000; // 9    **
		11'h69a: font_rom_data_out = 8'b00011000; // a    **
		11'h69b: font_rom_data_out = 8'b00111100; // b   ****
		11'h69c: font_rom_data_out = 8'b00000000; // c
		11'h69d: font_rom_data_out = 8'b00000000; // d
		11'h69e: font_rom_data_out = 8'b00000000; // e
		11'h69f: font_rom_data_out = 8'b00000000; // f
		// code x6a
		11'h6a0: font_rom_data_out = 8'b00000000; // 0
		11'h6a1: font_rom_data_out = 8'b00000000; // 1
		11'h6a2: font_rom_data_out = 8'b00000110; // 2      **
		11'h6a3: font_rom_data_out = 8'b00000110; // 3      **
		11'h6a4: font_rom_data_out = 8'b00000000; // 4
		11'h6a5: font_rom_data_out = 8'b00001110; // 5     ***
		11'h6a6: font_rom_data_out = 8'b00000110; // 6      **
		11'h6a7: font_rom_data_out = 8'b00000110; // 7      **
		11'h6a8: font_rom_data_out = 8'b00000110; // 8      **
		11'h6a9: font_rom_data_out = 8'b00000110; // 9      **
		11'h6aa: font_rom_data_out = 8'b00000110; // a      **
		11'h6ab: font_rom_data_out = 8'b00000110; // b      **
		11'h6ac: font_rom_data_out = 8'b01100110; // c  **  **
		11'h6ad: font_rom_data_out = 8'b01100110; // d  **  **
		11'h6ae: font_rom_data_out = 8'b00111100; // e   ****
		11'h6af: font_rom_data_out = 8'b00000000; // f
		// code x6b
		11'h6b0: font_rom_data_out = 8'b00000000; // 0
		11'h6b1: font_rom_data_out = 8'b00000000; // 1
		11'h6b2: font_rom_data_out = 8'b11100000; // 2 ***
		11'h6b3: font_rom_data_out = 8'b01100000; // 3  **
		11'h6b4: font_rom_data_out = 8'b01100000; // 4  **
		11'h6b5: font_rom_data_out = 8'b01100110; // 5  **  **
		11'h6b6: font_rom_data_out = 8'b01101100; // 6  ** **
		11'h6b7: font_rom_data_out = 8'b01111000; // 7  ****
		11'h6b8: font_rom_data_out = 8'b01111000; // 8  ****
		11'h6b9: font_rom_data_out = 8'b01101100; // 9  ** **
		11'h6ba: font_rom_data_out = 8'b01100110; // a  **  **
		11'h6bb: font_rom_data_out = 8'b11100110; // b ***  **
		11'h6bc: font_rom_data_out = 8'b00000000; // c
		11'h6bd: font_rom_data_out = 8'b00000000; // d
		11'h6be: font_rom_data_out = 8'b00000000; // e
		11'h6bf: font_rom_data_out = 8'b00000000; // f
		// code x6c
		11'h6c0: font_rom_data_out = 8'b00000000; // 0
		11'h6c1: font_rom_data_out = 8'b00000000; // 1
		11'h6c2: font_rom_data_out = 8'b00111000; // 2   ***
		11'h6c3: font_rom_data_out = 8'b00011000; // 3    **
		11'h6c4: font_rom_data_out = 8'b00011000; // 4    **
		11'h6c5: font_rom_data_out = 8'b00011000; // 5    **
		11'h6c6: font_rom_data_out = 8'b00011000; // 6    **
		11'h6c7: font_rom_data_out = 8'b00011000; // 7    **
		11'h6c8: font_rom_data_out = 8'b00011000; // 8    **
		11'h6c9: font_rom_data_out = 8'b00011000; // 9    **
		11'h6ca: font_rom_data_out = 8'b00011000; // a    **
		11'h6cb: font_rom_data_out = 8'b00111100; // b   ****
		11'h6cc: font_rom_data_out = 8'b00000000; // c
		11'h6cd: font_rom_data_out = 8'b00000000; // d
		11'h6ce: font_rom_data_out = 8'b00000000; // e
		11'h6cf: font_rom_data_out = 8'b00000000; // f
		// code x6d
		11'h6d0: font_rom_data_out = 8'b00000000; // 0
		11'h6d1: font_rom_data_out = 8'b00000000; // 1
		11'h6d2: font_rom_data_out = 8'b00000000; // 2
		11'h6d3: font_rom_data_out = 8'b00000000; // 3
		11'h6d4: font_rom_data_out = 8'b00000000; // 4
		11'h6d5: font_rom_data_out = 8'b11100110; // 5 ***  **
		11'h6d6: font_rom_data_out = 8'b11111111; // 6 ********
		11'h6d7: font_rom_data_out = 8'b11011011; // 7 ** ** **
		11'h6d8: font_rom_data_out = 8'b11011011; // 8 ** ** **
		11'h6d9: font_rom_data_out = 8'b11011011; // 9 ** ** **
		11'h6da: font_rom_data_out = 8'b11011011; // a ** ** **
		11'h6db: font_rom_data_out = 8'b11011011; // b ** ** **
		11'h6dc: font_rom_data_out = 8'b00000000; // c
		11'h6dd: font_rom_data_out = 8'b00000000; // d
		11'h6de: font_rom_data_out = 8'b00000000; // e
		11'h6df: font_rom_data_out = 8'b00000000; // f
		// code x6e
		11'h6e0: font_rom_data_out = 8'b00000000; // 0
		11'h6e1: font_rom_data_out = 8'b00000000; // 1
		11'h6e2: font_rom_data_out = 8'b00000000; // 2
		11'h6e3: font_rom_data_out = 8'b00000000; // 3
		11'h6e4: font_rom_data_out = 8'b00000000; // 4
		11'h6e5: font_rom_data_out = 8'b11011100; // 5 ** ***
		11'h6e6: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h6e7: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h6e8: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h6e9: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h6ea: font_rom_data_out = 8'b01100110; // a  **  **
		11'h6eb: font_rom_data_out = 8'b01100110; // b  **  **
		11'h6ec: font_rom_data_out = 8'b00000000; // c
		11'h6ed: font_rom_data_out = 8'b00000000; // d
		11'h6ee: font_rom_data_out = 8'b00000000; // e
		11'h6ef: font_rom_data_out = 8'b00000000; // f
		// code x6f
		11'h6f0: font_rom_data_out = 8'b00000000; // 0
		11'h6f1: font_rom_data_out = 8'b00000000; // 1
		11'h6f2: font_rom_data_out = 8'b00000000; // 2
		11'h6f3: font_rom_data_out = 8'b00000000; // 3
		11'h6f4: font_rom_data_out = 8'b00000000; // 4
		11'h6f5: font_rom_data_out = 8'b01111100; // 5  *****
		11'h6f6: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h6f7: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h6f8: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h6f9: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h6fa: font_rom_data_out = 8'b11000110; // a **   **
		11'h6fb: font_rom_data_out = 8'b01111100; // b  *****
		11'h6fc: font_rom_data_out = 8'b00000000; // c
		11'h6fd: font_rom_data_out = 8'b00000000; // d
		11'h6fe: font_rom_data_out = 8'b00000000; // e
		11'h6ff: font_rom_data_out = 8'b00000000; // f
		// code x70
		11'h700: font_rom_data_out = 8'b00000000; // 0
		11'h701: font_rom_data_out = 8'b00000000; // 1
		11'h702: font_rom_data_out = 8'b00000000; // 2
		11'h703: font_rom_data_out = 8'b00000000; // 3
		11'h704: font_rom_data_out = 8'b00000000; // 4
		11'h705: font_rom_data_out = 8'b11011100; // 5 ** ***
		11'h706: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h707: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h708: font_rom_data_out = 8'b01100110; // 8  **  **
		11'h709: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h70a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h70b: font_rom_data_out = 8'b01111100; // b  *****
		11'h70c: font_rom_data_out = 8'b01100000; // c  **
		11'h70d: font_rom_data_out = 8'b01100000; // d  **
		11'h70e: font_rom_data_out = 8'b11110000; // e ****
		11'h70f: font_rom_data_out = 8'b00000000; // f
		// code x71
		11'h710: font_rom_data_out = 8'b00000000; // 0
		11'h711: font_rom_data_out = 8'b00000000; // 1
		11'h712: font_rom_data_out = 8'b00000000; // 2
		11'h713: font_rom_data_out = 8'b00000000; // 3
		11'h714: font_rom_data_out = 8'b00000000; // 4
		11'h715: font_rom_data_out = 8'b01110110; // 5  *** **
		11'h716: font_rom_data_out = 8'b11001100; // 6 **  **
		11'h717: font_rom_data_out = 8'b11001100; // 7 **  **
		11'h718: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h719: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h71a: font_rom_data_out = 8'b11001100; // a **  **
		11'h71b: font_rom_data_out = 8'b01111100; // b  *****
		11'h71c: font_rom_data_out = 8'b00001100; // c     **
		11'h71d: font_rom_data_out = 8'b00001100; // d     **
		11'h71e: font_rom_data_out = 8'b00011110; // e    ****
		11'h71f: font_rom_data_out = 8'b00000000; // f
		// code x72
		11'h720: font_rom_data_out = 8'b00000000; // 0
		11'h721: font_rom_data_out = 8'b00000000; // 1
		11'h722: font_rom_data_out = 8'b00000000; // 2
		11'h723: font_rom_data_out = 8'b00000000; // 3
		11'h724: font_rom_data_out = 8'b00000000; // 4
		11'h725: font_rom_data_out = 8'b11011100; // 5 ** ***
		11'h726: font_rom_data_out = 8'b01110110; // 6  *** **
		11'h727: font_rom_data_out = 8'b01100110; // 7  **  **
		11'h728: font_rom_data_out = 8'b01100000; // 8  **
		11'h729: font_rom_data_out = 8'b01100000; // 9  **
		11'h72a: font_rom_data_out = 8'b01100000; // a  **
		11'h72b: font_rom_data_out = 8'b11110000; // b ****
		11'h72c: font_rom_data_out = 8'b00000000; // c
		11'h72d: font_rom_data_out = 8'b00000000; // d
		11'h72e: font_rom_data_out = 8'b00000000; // e
		11'h72f: font_rom_data_out = 8'b00000000; // f
		// code x73
		11'h730: font_rom_data_out = 8'b00000000; // 0
		11'h731: font_rom_data_out = 8'b00000000; // 1
		11'h732: font_rom_data_out = 8'b00000000; // 2
		11'h733: font_rom_data_out = 8'b00000000; // 3
		11'h734: font_rom_data_out = 8'b00000000; // 4
		11'h735: font_rom_data_out = 8'b01111100; // 5  *****
		11'h736: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h737: font_rom_data_out = 8'b01100000; // 7  **
		11'h738: font_rom_data_out = 8'b00111000; // 8   ***
		11'h739: font_rom_data_out = 8'b00001100; // 9     **
		11'h73a: font_rom_data_out = 8'b11000110; // a **   **
		11'h73b: font_rom_data_out = 8'b01111100; // b  *****
		11'h73c: font_rom_data_out = 8'b00000000; // c
		11'h73d: font_rom_data_out = 8'b00000000; // d
		11'h73e: font_rom_data_out = 8'b00000000; // e
		11'h73f: font_rom_data_out = 8'b00000000; // f
		// code x74
		11'h740: font_rom_data_out = 8'b00000000; // 0
		11'h741: font_rom_data_out = 8'b00000000; // 1
		11'h742: font_rom_data_out = 8'b00010000; // 2    *
		11'h743: font_rom_data_out = 8'b00110000; // 3   **
		11'h744: font_rom_data_out = 8'b00110000; // 4   **
		11'h745: font_rom_data_out = 8'b11111100; // 5 ******
		11'h746: font_rom_data_out = 8'b00110000; // 6   **
		11'h747: font_rom_data_out = 8'b00110000; // 7   **
		11'h748: font_rom_data_out = 8'b00110000; // 8   **
		11'h749: font_rom_data_out = 8'b00110000; // 9   **
		11'h74a: font_rom_data_out = 8'b00110110; // a   ** **
		11'h74b: font_rom_data_out = 8'b00011100; // b    ***
		11'h74c: font_rom_data_out = 8'b00000000; // c
		11'h74d: font_rom_data_out = 8'b00000000; // d
		11'h74e: font_rom_data_out = 8'b00000000; // e
		11'h74f: font_rom_data_out = 8'b00000000; // f
		// code x75
		11'h750: font_rom_data_out = 8'b00000000; // 0
		11'h751: font_rom_data_out = 8'b00000000; // 1
		11'h752: font_rom_data_out = 8'b00000000; // 2
		11'h753: font_rom_data_out = 8'b00000000; // 3
		11'h754: font_rom_data_out = 8'b00000000; // 4
		11'h755: font_rom_data_out = 8'b11001100; // 5 **  **
		11'h756: font_rom_data_out = 8'b11001100; // 6 **  **
		11'h757: font_rom_data_out = 8'b11001100; // 7 **  **
		11'h758: font_rom_data_out = 8'b11001100; // 8 **  **
		11'h759: font_rom_data_out = 8'b11001100; // 9 **  **
		11'h75a: font_rom_data_out = 8'b11001100; // a **  **
		11'h75b: font_rom_data_out = 8'b01110110; // b  *** **
		11'h75c: font_rom_data_out = 8'b00000000; // c
		11'h75d: font_rom_data_out = 8'b00000000; // d
		11'h75e: font_rom_data_out = 8'b00000000; // e
		11'h75f: font_rom_data_out = 8'b00000000; // f
		// code x76
		11'h760: font_rom_data_out = 8'b00000000; // 0
		11'h761: font_rom_data_out = 8'b00000000; // 1
		11'h762: font_rom_data_out = 8'b00000000; // 2
		11'h763: font_rom_data_out = 8'b00000000; // 3
		11'h764: font_rom_data_out = 8'b00000000; // 4
		11'h765: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h766: font_rom_data_out = 8'b11000011; // 6 **    **
		11'h767: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h768: font_rom_data_out = 8'b11000011; // 8 **    **
		11'h769: font_rom_data_out = 8'b01100110; // 9  **  **
		11'h76a: font_rom_data_out = 8'b00111100; // a   ****
		11'h76b: font_rom_data_out = 8'b00011000; // b    **
		11'h76c: font_rom_data_out = 8'b00000000; // c
		11'h76d: font_rom_data_out = 8'b00000000; // d
		11'h76e: font_rom_data_out = 8'b00000000; // e
		11'h76f: font_rom_data_out = 8'b00000000; // f
		// code x77
		11'h770: font_rom_data_out = 8'b00000000; // 0
		11'h771: font_rom_data_out = 8'b00000000; // 1
		11'h772: font_rom_data_out = 8'b00000000; // 2
		11'h773: font_rom_data_out = 8'b00000000; // 3
		11'h774: font_rom_data_out = 8'b00000000; // 4
		11'h775: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h776: font_rom_data_out = 8'b11000011; // 6 **    **
		11'h777: font_rom_data_out = 8'b11000011; // 7 **    **
		11'h778: font_rom_data_out = 8'b11011011; // 8 ** ** **
		11'h779: font_rom_data_out = 8'b11011011; // 9 ** ** **
		11'h77a: font_rom_data_out = 8'b11111111; // a ********
		11'h77b: font_rom_data_out = 8'b01100110; // b  **  **
		11'h77c: font_rom_data_out = 8'b00000000; // c
		11'h77d: font_rom_data_out = 8'b00000000; // d
		11'h77e: font_rom_data_out = 8'b00000000; // e
		11'h77f: font_rom_data_out = 8'b00000000; // f
		// code x78
		11'h780: font_rom_data_out = 8'b00000000; // 0
		11'h781: font_rom_data_out = 8'b00000000; // 1
		11'h782: font_rom_data_out = 8'b00000000; // 2
		11'h783: font_rom_data_out = 8'b00000000; // 3
		11'h784: font_rom_data_out = 8'b00000000; // 4
		11'h785: font_rom_data_out = 8'b11000011; // 5 **    **
		11'h786: font_rom_data_out = 8'b01100110; // 6  **  **
		11'h787: font_rom_data_out = 8'b00111100; // 7   ****
		11'h788: font_rom_data_out = 8'b00011000; // 8    **
		11'h789: font_rom_data_out = 8'b00111100; // 9   ****
		11'h78a: font_rom_data_out = 8'b01100110; // a  **  **
		11'h78b: font_rom_data_out = 8'b11000011; // b **    **
		11'h78c: font_rom_data_out = 8'b00000000; // c
		11'h78d: font_rom_data_out = 8'b00000000; // d
		11'h78e: font_rom_data_out = 8'b00000000; // e
		11'h78f: font_rom_data_out = 8'b00000000; // f
		// code x79
		11'h790: font_rom_data_out = 8'b00000000; // 0
		11'h791: font_rom_data_out = 8'b00000000; // 1
		11'h792: font_rom_data_out = 8'b00000000; // 2
		11'h793: font_rom_data_out = 8'b00000000; // 3
		11'h794: font_rom_data_out = 8'b00000000; // 4
		11'h795: font_rom_data_out = 8'b11000110; // 5 **   **
		11'h796: font_rom_data_out = 8'b11000110; // 6 **   **
		11'h797: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h798: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h799: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h79a: font_rom_data_out = 8'b11000110; // a **   **
		11'h79b: font_rom_data_out = 8'b01111110; // b  ******
		11'h79c: font_rom_data_out = 8'b00000110; // c      **
		11'h79d: font_rom_data_out = 8'b00001100; // d     **
		11'h79e: font_rom_data_out = 8'b11111000; // e *****
		11'h79f: font_rom_data_out = 8'b00000000; // f
		// code x7a
		11'h7a0: font_rom_data_out = 8'b00000000; // 0
		11'h7a1: font_rom_data_out = 8'b00000000; // 1
		11'h7a2: font_rom_data_out = 8'b00000000; // 2
		11'h7a3: font_rom_data_out = 8'b00000000; // 3
		11'h7a4: font_rom_data_out = 8'b00000000; // 4
		11'h7a5: font_rom_data_out = 8'b11111110; // 5 *******
		11'h7a6: font_rom_data_out = 8'b11001100; // 6 **  **
		11'h7a7: font_rom_data_out = 8'b00011000; // 7    **
		11'h7a8: font_rom_data_out = 8'b00110000; // 8   **
		11'h7a9: font_rom_data_out = 8'b01100000; // 9  **
		11'h7aa: font_rom_data_out = 8'b11000110; // a **   **
		11'h7ab: font_rom_data_out = 8'b11111110; // b *******
		11'h7ac: font_rom_data_out = 8'b00000000; // c
		11'h7ad: font_rom_data_out = 8'b00000000; // d
		11'h7ae: font_rom_data_out = 8'b00000000; // e
		11'h7af: font_rom_data_out = 8'b00000000; // f
		// code x7b
		11'h7b0: font_rom_data_out = 8'b00000000; // 0
		11'h7b1: font_rom_data_out = 8'b00000000; // 1
		11'h7b2: font_rom_data_out = 8'b00001110; // 2     ***
		11'h7b3: font_rom_data_out = 8'b00011000; // 3    **
		11'h7b4: font_rom_data_out = 8'b00011000; // 4    **
		11'h7b5: font_rom_data_out = 8'b00011000; // 5    **
		11'h7b6: font_rom_data_out = 8'b01110000; // 6  ***
		11'h7b7: font_rom_data_out = 8'b00011000; // 7    **
		11'h7b8: font_rom_data_out = 8'b00011000; // 8    **
		11'h7b9: font_rom_data_out = 8'b00011000; // 9    **
		11'h7ba: font_rom_data_out = 8'b00011000; // a    **
		11'h7bb: font_rom_data_out = 8'b00001110; // b     ***
		11'h7bc: font_rom_data_out = 8'b00000000; // c
		11'h7bd: font_rom_data_out = 8'b00000000; // d
		11'h7be: font_rom_data_out = 8'b00000000; // e
		11'h7bf: font_rom_data_out = 8'b00000000; // f
		// code x7c
		11'h7c0: font_rom_data_out = 8'b00000000; // 0
		11'h7c1: font_rom_data_out = 8'b00000000; // 1
		11'h7c2: font_rom_data_out = 8'b00011000; // 2    **
		11'h7c3: font_rom_data_out = 8'b00011000; // 3    **
		11'h7c4: font_rom_data_out = 8'b00011000; // 4    **
		11'h7c5: font_rom_data_out = 8'b00011000; // 5    **
		11'h7c6: font_rom_data_out = 8'b00000000; // 6
		11'h7c7: font_rom_data_out = 8'b00011000; // 7    **
		11'h7c8: font_rom_data_out = 8'b00011000; // 8    **
		11'h7c9: font_rom_data_out = 8'b00011000; // 9    **
		11'h7ca: font_rom_data_out = 8'b00011000; // a    **
		11'h7cb: font_rom_data_out = 8'b00011000; // b    **
		11'h7cc: font_rom_data_out = 8'b00000000; // c
		11'h7cd: font_rom_data_out = 8'b00000000; // d
		11'h7ce: font_rom_data_out = 8'b00000000; // e
		11'h7cf: font_rom_data_out = 8'b00000000; // f
		// code x7d
		11'h7d0: font_rom_data_out = 8'b00000000; // 0
		11'h7d1: font_rom_data_out = 8'b00000000; // 1
		11'h7d2: font_rom_data_out = 8'b01110000; // 2  ***
		11'h7d3: font_rom_data_out = 8'b00011000; // 3    **
		11'h7d4: font_rom_data_out = 8'b00011000; // 4    **
		11'h7d5: font_rom_data_out = 8'b00011000; // 5    **
		11'h7d6: font_rom_data_out = 8'b00001110; // 6     ***
		11'h7d7: font_rom_data_out = 8'b00011000; // 7    **
		11'h7d8: font_rom_data_out = 8'b00011000; // 8    **
		11'h7d9: font_rom_data_out = 8'b00011000; // 9    **
		11'h7da: font_rom_data_out = 8'b00011000; // a    **
		11'h7db: font_rom_data_out = 8'b01110000; // b  ***
		11'h7dc: font_rom_data_out = 8'b00000000; // c
		11'h7dd: font_rom_data_out = 8'b00000000; // d
		11'h7de: font_rom_data_out = 8'b00000000; // e
		11'h7df: font_rom_data_out = 8'b00000000; // f
		// code x7e
		11'h7e0: font_rom_data_out = 8'b00000000; // 0
		11'h7e1: font_rom_data_out = 8'b00000000; // 1
		11'h7e2: font_rom_data_out = 8'b01110110; // 2  *** **
		11'h7e3: font_rom_data_out = 8'b11011100; // 3 ** ***
		11'h7e4: font_rom_data_out = 8'b00000000; // 4
		11'h7e5: font_rom_data_out = 8'b00000000; // 5
		11'h7e6: font_rom_data_out = 8'b00000000; // 6
		11'h7e7: font_rom_data_out = 8'b00000000; // 7
		11'h7e8: font_rom_data_out = 8'b00000000; // 8
		11'h7e9: font_rom_data_out = 8'b00000000; // 9
		11'h7ea: font_rom_data_out = 8'b00000000; // a
		11'h7eb: font_rom_data_out = 8'b00000000; // b
		11'h7ec: font_rom_data_out = 8'b00000000; // c
		11'h7ed: font_rom_data_out = 8'b00000000; // d
		11'h7ee: font_rom_data_out = 8'b00000000; // e
		11'h7ef: font_rom_data_out = 8'b00000000; // f
		// code x7f
		11'h7f0: font_rom_data_out = 8'b00000000; // 0
		11'h7f1: font_rom_data_out = 8'b00000000; // 1
		11'h7f2: font_rom_data_out = 8'b00000000; // 2
		11'h7f3: font_rom_data_out = 8'b00000000; // 3
		11'h7f4: font_rom_data_out = 8'b00010000; // 4    *
		11'h7f5: font_rom_data_out = 8'b00111000; // 5   ***
		11'h7f6: font_rom_data_out = 8'b01101100; // 6  ** **
		11'h7f7: font_rom_data_out = 8'b11000110; // 7 **   **
		11'h7f8: font_rom_data_out = 8'b11000110; // 8 **   **
		11'h7f9: font_rom_data_out = 8'b11000110; // 9 **   **
		11'h7fa: font_rom_data_out = 8'b11111110; // a *******
		11'h7fb: font_rom_data_out = 8'b00000000; // b
		11'h7fc: font_rom_data_out = 8'b00000000; // c
		11'h7fd: font_rom_data_out = 8'b00000000; // d
		11'h7fe: font_rom_data_out = 8'b00000000; // e
		11'h7ff: font_rom_data_out = 8'b00000000; // f
        default: font_rom_data_out = 8'b00000000;
    endcase
endmodule