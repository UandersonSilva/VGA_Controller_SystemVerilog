module  font_rom ( 
        //input logic font_rom_clk_in,  
        input logic [10:0] addr_in,  
        output logic [7:0] data_out
    ); 
  
    //logic [10:0] addr_reg;

    //always_ff @(posedge font_rom_clk_in)
	always @(addr_in)
	begin
       //addr_reg <= addr_in;

		case(addr_in)
			11'h000: data_out = 8'b00000000; // 0
			11'h001: data_out = 8'b00000000; // 1
			11'h002: data_out = 8'b00000000; // 2
			11'h003: data_out = 8'b00000000; // 3
			11'h004: data_out = 8'b00000000; // 4
			11'h005: data_out = 8'b00000000; // 5
			11'h006: data_out = 8'b00000000; // 6
			11'h007: data_out = 8'b00000000; // 7
			11'h008: data_out = 8'b00000000; // 8
			11'h009: data_out = 8'b00000000; // 9
			11'h00a: data_out = 8'b00000000; // a
			11'h00b: data_out = 8'b00000000; // b
			11'h00c: data_out = 8'b00000000; // c
			11'h00d: data_out = 8'b00000000; // d
			11'h00e: data_out = 8'b00000000; // e
			11'h00f: data_out = 8'b00000000; // f
			// code x01
			11'h010: data_out = 8'b00000000; // 0
			11'h011: data_out = 8'b00000000; // 1
			11'h012: data_out = 8'b01111110; // 2  ******
			11'h013: data_out = 8'b10000001; // 3 *      *
			11'h014: data_out = 8'b10100101; // 4 * *  * *
			11'h015: data_out = 8'b10000001; // 5 *      *
			11'h016: data_out = 8'b10000001; // 6 *      *
			11'h017: data_out = 8'b10111101; // 7 * **** *
			11'h018: data_out = 8'b10011001; // 8 *  **  *
			11'h019: data_out = 8'b10000001; // 9 *      *
			11'h01a: data_out = 8'b10000001; // a *      *
			11'h01b: data_out = 8'b01111110; // b  ******
			11'h01c: data_out = 8'b00000000; // c
			11'h01d: data_out = 8'b00000000; // d
			11'h01e: data_out = 8'b00000000; // e
			11'h01f: data_out = 8'b00000000; // f
			// code x02
			11'h020: data_out = 8'b00000000; // 0
			11'h021: data_out = 8'b00000000; // 1
			11'h022: data_out = 8'b01111110; // 2  ******
			11'h023: data_out = 8'b11111111; // 3 ********
			11'h024: data_out = 8'b11011011; // 4 ** ** **
			11'h025: data_out = 8'b11111111; // 5 ********
			11'h026: data_out = 8'b11111111; // 6 ********
			11'h027: data_out = 8'b11000011; // 7 **    **
			11'h028: data_out = 8'b11100111; // 8 ***  ***
			11'h029: data_out = 8'b11111111; // 9 ********
			11'h02a: data_out = 8'b11111111; // a ********
			11'h02b: data_out = 8'b01111110; // b  ******
			11'h02c: data_out = 8'b00000000; // c
			11'h02d: data_out = 8'b00000000; // d
			11'h02e: data_out = 8'b00000000; // e
			11'h02f: data_out = 8'b00000000; // f
			// code x03
			11'h030: data_out = 8'b00000000; // 0
			11'h031: data_out = 8'b00000000; // 1
			11'h032: data_out = 8'b00000000; // 2
			11'h033: data_out = 8'b00000000; // 3
			11'h034: data_out = 8'b01101100; // 4  ** **
			11'h035: data_out = 8'b11111110; // 5 *******
			11'h036: data_out = 8'b11111110; // 6 *******
			11'h037: data_out = 8'b11111110; // 7 *******
			11'h038: data_out = 8'b11111110; // 8 *******
			11'h039: data_out = 8'b01111100; // 9  *****
			11'h03a: data_out = 8'b00111000; // a   ***
			11'h03b: data_out = 8'b00010000; // b    *
			11'h03c: data_out = 8'b00000000; // c
			11'h03d: data_out = 8'b00000000; // d
			11'h03e: data_out = 8'b00000000; // e
			11'h03f: data_out = 8'b00000000; // f
			// code x04
			11'h040: data_out = 8'b00000000; // 0
			11'h041: data_out = 8'b00000000; // 1
			11'h042: data_out = 8'b00000000; // 2
			11'h043: data_out = 8'b00000000; // 3
			11'h044: data_out = 8'b00010000; // 4    *
			11'h045: data_out = 8'b00111000; // 5   ***
			11'h046: data_out = 8'b01111100; // 6  *****
			11'h047: data_out = 8'b11111110; // 7 *******
			11'h048: data_out = 8'b01111100; // 8  *****
			11'h049: data_out = 8'b00111000; // 9   ***
			11'h04a: data_out = 8'b00010000; // a    *
			11'h04b: data_out = 8'b00000000; // b
			11'h04c: data_out = 8'b00000000; // c
			11'h04d: data_out = 8'b00000000; // d
			11'h04e: data_out = 8'b00000000; // e
			11'h04f: data_out = 8'b00000000; // f
			// code x05
			11'h050: data_out = 8'b00000000; // 0
			11'h051: data_out = 8'b00000000; // 1
			11'h052: data_out = 8'b00000000; // 2
			11'h053: data_out = 8'b00011000; // 3    **
			11'h054: data_out = 8'b00111100; // 4   ****
			11'h055: data_out = 8'b00111100; // 5   ****
			11'h056: data_out = 8'b11100111; // 6 ***  ***
			11'h057: data_out = 8'b11100111; // 7 ***  ***
			11'h058: data_out = 8'b11100111; // 8 ***  ***
			11'h059: data_out = 8'b00011000; // 9    **
			11'h05a: data_out = 8'b00011000; // a    **
			11'h05b: data_out = 8'b00111100; // b   ****
			11'h05c: data_out = 8'b00000000; // c
			11'h05d: data_out = 8'b00000000; // d
			11'h05e: data_out = 8'b00000000; // e
			11'h05f: data_out = 8'b00000000; // f
			// code x06
			11'h060: data_out = 8'b00000000; // 0
			11'h061: data_out = 8'b00000000; // 1
			11'h062: data_out = 8'b00000000; // 2
			11'h063: data_out = 8'b00011000; // 3    **
			11'h064: data_out = 8'b00111100; // 4   ****
			11'h065: data_out = 8'b01111110; // 5  ******
			11'h066: data_out = 8'b11111111; // 6 ********
			11'h067: data_out = 8'b11111111; // 7 ********
			11'h068: data_out = 8'b01111110; // 8  ******
			11'h069: data_out = 8'b00011000; // 9    **
			11'h06a: data_out = 8'b00011000; // a    **
			11'h06b: data_out = 8'b00111100; // b   ****
			11'h06c: data_out = 8'b00000000; // c
			11'h06d: data_out = 8'b00000000; // d
			11'h06e: data_out = 8'b00000000; // e
			11'h06f: data_out = 8'b00000000; // f
			// code x07
			11'h070: data_out = 8'b00000000; // 0
			11'h071: data_out = 8'b00000000; // 1
			11'h072: data_out = 8'b00000000; // 2
			11'h073: data_out = 8'b00000000; // 3
			11'h074: data_out = 8'b00000000; // 4
			11'h075: data_out = 8'b00000000; // 5
			11'h076: data_out = 8'b00011000; // 6    **
			11'h077: data_out = 8'b00111100; // 7   ****
			11'h078: data_out = 8'b00111100; // 8   ****
			11'h079: data_out = 8'b00011000; // 9    **
			11'h07a: data_out = 8'b00000000; // a
			11'h07b: data_out = 8'b00000000; // b
			11'h07c: data_out = 8'b00000000; // c
			11'h07d: data_out = 8'b00000000; // d
			11'h07e: data_out = 8'b00000000; // e
			11'h07f: data_out = 8'b00000000; // f
			// code x08
			11'h080: data_out = 8'b11111111; // 0 ********
			11'h081: data_out = 8'b11111111; // 1 ********
			11'h082: data_out = 8'b11111111; // 2 ********
			11'h083: data_out = 8'b11111111; // 3 ********
			11'h084: data_out = 8'b11111111; // 4 ********
			11'h085: data_out = 8'b11111111; // 5 ********
			11'h086: data_out = 8'b11100111; // 6 ***  ***
			11'h087: data_out = 8'b11000011; // 7 **    **
			11'h088: data_out = 8'b11000011; // 8 **    **
			11'h089: data_out = 8'b11100111; // 9 ***  ***
			11'h08a: data_out = 8'b11111111; // a ********
			11'h08b: data_out = 8'b11111111; // b ********
			11'h08c: data_out = 8'b11111111; // c ********
			11'h08d: data_out = 8'b11111111; // d ********
			11'h08e: data_out = 8'b11111111; // e ********
			11'h08f: data_out = 8'b11111111; // f ********
			// code x09
			11'h090: data_out = 8'b00000000; // 0
			11'h091: data_out = 8'b00000000; // 1
			11'h092: data_out = 8'b00000000; // 2
			11'h093: data_out = 8'b00000000; // 3
			11'h094: data_out = 8'b00000000; // 4
			11'h095: data_out = 8'b00111100; // 5   ****
			11'h096: data_out = 8'b01100110; // 6  **  **
			11'h097: data_out = 8'b01000010; // 7  *    *
			11'h098: data_out = 8'b01000010; // 8  *    *
			11'h099: data_out = 8'b01100110; // 9  **  **
			11'h09a: data_out = 8'b00111100; // a   ****
			11'h09b: data_out = 8'b00000000; // b
			11'h09c: data_out = 8'b00000000; // c
			11'h09d: data_out = 8'b00000000; // d
			11'h09e: data_out = 8'b00000000; // e
			11'h09f: data_out = 8'b00000000; // f
			// code x0a
			11'h0a0: data_out = 8'b11111111; // 0 ********
			11'h0a1: data_out = 8'b11111111; // 1 ********
			11'h0a2: data_out = 8'b11111111; // 2 ********
			11'h0a3: data_out = 8'b11111111; // 3 ********
			11'h0a4: data_out = 8'b11111111; // 4 ********
			11'h0a5: data_out = 8'b11000011; // 5 **    **
			11'h0a6: data_out = 8'b10011001; // 6 *  **  *
			11'h0a7: data_out = 8'b10111101; // 7 * **** *
			11'h0a8: data_out = 8'b10111101; // 8 * **** *
			11'h0a9: data_out = 8'b10011001; // 9 *  **  *
			11'h0aa: data_out = 8'b11000011; // a **    **
			11'h0ab: data_out = 8'b11111111; // b ********
			11'h0ac: data_out = 8'b11111111; // c ********
			11'h0ad: data_out = 8'b11111111; // d ********
			11'h0ae: data_out = 8'b11111111; // e ********
			11'h0af: data_out = 8'b11111111; // f ********
			// code x0b
			11'h0b0: data_out = 8'b00000000; // 0
			11'h0b1: data_out = 8'b00000000; // 1
			11'h0b2: data_out = 8'b00011110; // 2    ****
			11'h0b3: data_out = 8'b00001110; // 3     ***
			11'h0b4: data_out = 8'b00011010; // 4    ** *
			11'h0b5: data_out = 8'b00110010; // 5   **  *
			11'h0b6: data_out = 8'b01111000; // 6  ****
			11'h0b7: data_out = 8'b11001100; // 7 **  **
			11'h0b8: data_out = 8'b11001100; // 8 **  **
			11'h0b9: data_out = 8'b11001100; // 9 **  **
			11'h0ba: data_out = 8'b11001100; // a **  **
			11'h0bb: data_out = 8'b01111000; // b  ****
			11'h0bc: data_out = 8'b00000000; // c
			11'h0bd: data_out = 8'b00000000; // d
			11'h0be: data_out = 8'b00000000; // e
			11'h0bf: data_out = 8'b00000000; // f
			// code x0c
			11'h0c0: data_out = 8'b00000000; // 0
			11'h0c1: data_out = 8'b00000000; // 1
			11'h0c2: data_out = 8'b00111100; // 2   ****
			11'h0c3: data_out = 8'b01100110; // 3  **  **
			11'h0c4: data_out = 8'b01100110; // 4  **  **
			11'h0c5: data_out = 8'b01100110; // 5  **  **
			11'h0c6: data_out = 8'b01100110; // 6  **  **
			11'h0c7: data_out = 8'b00111100; // 7   ****
			11'h0c8: data_out = 8'b00011000; // 8    **
			11'h0c9: data_out = 8'b01111110; // 9  ******
			11'h0ca: data_out = 8'b00011000; // a    **
			11'h0cb: data_out = 8'b00011000; // b    **
			11'h0cc: data_out = 8'b00000000; // c
			11'h0cd: data_out = 8'b00000000; // d
			11'h0ce: data_out = 8'b00000000; // e
			11'h0cf: data_out = 8'b00000000; // f
			// code x0d
			11'h0d0: data_out = 8'b00000000; // 0
			11'h0d1: data_out = 8'b00000000; // 1
			11'h0d2: data_out = 8'b00111111; // 2   ******
			11'h0d3: data_out = 8'b00110011; // 3   **  **
			11'h0d4: data_out = 8'b00111111; // 4   ******
			11'h0d5: data_out = 8'b00110000; // 5   **
			11'h0d6: data_out = 8'b00110000; // 6   **
			11'h0d7: data_out = 8'b00110000; // 7   **
			11'h0d8: data_out = 8'b00110000; // 8   **
			11'h0d9: data_out = 8'b01110000; // 9  ***
			11'h0da: data_out = 8'b11110000; // a ****
			11'h0db: data_out = 8'b11100000; // b ***
			11'h0dc: data_out = 8'b00000000; // c
			11'h0dd: data_out = 8'b00000000; // d
			11'h0de: data_out = 8'b00000000; // e
			11'h0df: data_out = 8'b00000000; // f
			// code x0e
			11'h0e0: data_out = 8'b00000000; // 0
			11'h0e1: data_out = 8'b00000000; // 1
			11'h0e2: data_out = 8'b01111111; // 2  *******
			11'h0e3: data_out = 8'b01100011; // 3  **   **
			11'h0e4: data_out = 8'b01111111; // 4  *******
			11'h0e5: data_out = 8'b01100011; // 5  **   **
			11'h0e6: data_out = 8'b01100011; // 6  **   **
			11'h0e7: data_out = 8'b01100011; // 7  **   **
			11'h0e8: data_out = 8'b01100011; // 8  **   **
			11'h0e9: data_out = 8'b01100111; // 9  **  ***
			11'h0ea: data_out = 8'b11100111; // a ***  ***
			11'h0eb: data_out = 8'b11100110; // b ***  **
			11'h0ec: data_out = 8'b11000000; // c **
			11'h0ed: data_out = 8'b00000000; // d
			11'h0ee: data_out = 8'b00000000; // e
			11'h0ef: data_out = 8'b00000000; // f
			// code x0f
			11'h0f0: data_out = 8'b00000000; // 0
			11'h0f1: data_out = 8'b00000000; // 1
			11'h0f2: data_out = 8'b00000000; // 2
			11'h0f3: data_out = 8'b00011000; // 3    **
			11'h0f4: data_out = 8'b00011000; // 4    **
			11'h0f5: data_out = 8'b11011011; // 5 ** ** **
			11'h0f6: data_out = 8'b00111100; // 6   ****
			11'h0f7: data_out = 8'b11100111; // 7 ***  ***
			11'h0f8: data_out = 8'b00111100; // 8   ****
			11'h0f9: data_out = 8'b11011011; // 9 ** ** **
			11'h0fa: data_out = 8'b00011000; // a    **
			11'h0fb: data_out = 8'b00011000; // b    **
			11'h0fc: data_out = 8'b00000000; // c
			11'h0fd: data_out = 8'b00000000; // d
			11'h0fe: data_out = 8'b00000000; // e
			11'h0ff: data_out = 8'b00000000; // f
			// code x10
			11'h100: data_out = 8'b00000000; // 0
			11'h101: data_out = 8'b10000000; // 1 *
			11'h102: data_out = 8'b11000000; // 2 **
			11'h103: data_out = 8'b11100000; // 3 ***
			11'h104: data_out = 8'b11110000; // 4 ****
			11'h105: data_out = 8'b11111000; // 5 *****
			11'h106: data_out = 8'b11111110; // 6 *******
			11'h107: data_out = 8'b11111000; // 7 *****
			11'h108: data_out = 8'b11110000; // 8 ****
			11'h109: data_out = 8'b11100000; // 9 ***
			11'h10a: data_out = 8'b11000000; // a **
			11'h10b: data_out = 8'b10000000; // b *
			11'h10c: data_out = 8'b00000000; // c
			11'h10d: data_out = 8'b00000000; // d
			11'h10e: data_out = 8'b00000000; // e
			11'h10f: data_out = 8'b00000000; // f
			// code x11
			11'h110: data_out = 8'b00000000; // 0
			11'h111: data_out = 8'b00000010; // 1       *
			11'h112: data_out = 8'b00000110; // 2      **
			11'h113: data_out = 8'b00001110; // 3     ***
			11'h114: data_out = 8'b00011110; // 4    ****
			11'h115: data_out = 8'b00111110; // 5   *****
			11'h116: data_out = 8'b11111110; // 6 *******
			11'h117: data_out = 8'b00111110; // 7   *****
			11'h118: data_out = 8'b00011110; // 8    ****
			11'h119: data_out = 8'b00001110; // 9     ***
			11'h11a: data_out = 8'b00000110; // a      **
			11'h11b: data_out = 8'b00000010; // b       *
			11'h11c: data_out = 8'b00000000; // c
			11'h11d: data_out = 8'b00000000; // d
			11'h11e: data_out = 8'b00000000; // e
			11'h11f: data_out = 8'b00000000; // f
			// code x12
			11'h120: data_out = 8'b00000000; // 0
			11'h121: data_out = 8'b00000000; // 1
			11'h122: data_out = 8'b00011000; // 2    **
			11'h123: data_out = 8'b00111100; // 3   ****
			11'h124: data_out = 8'b01111110; // 4  ******
			11'h125: data_out = 8'b00011000; // 5    **
			11'h126: data_out = 8'b00011000; // 6    **
			11'h127: data_out = 8'b00011000; // 7    **
			11'h128: data_out = 8'b01111110; // 8  ******
			11'h129: data_out = 8'b00111100; // 9   ****
			11'h12a: data_out = 8'b00011000; // a    **
			11'h12b: data_out = 8'b00000000; // b
			11'h12c: data_out = 8'b00000000; // c
			11'h12d: data_out = 8'b00000000; // d
			11'h12e: data_out = 8'b00000000; // e
			11'h12f: data_out = 8'b00000000; // f
			// code x13
			11'h130: data_out = 8'b00000000; // 0
			11'h131: data_out = 8'b00000000; // 1
			11'h132: data_out = 8'b01100110; // 2  **  **
			11'h133: data_out = 8'b01100110; // 3  **  **
			11'h134: data_out = 8'b01100110; // 4  **  **
			11'h135: data_out = 8'b01100110; // 5  **  **
			11'h136: data_out = 8'b01100110; // 6  **  **
			11'h137: data_out = 8'b01100110; // 7  **  **
			11'h138: data_out = 8'b01100110; // 8  **  **
			11'h139: data_out = 8'b00000000; // 9
			11'h13a: data_out = 8'b01100110; // a  **  **
			11'h13b: data_out = 8'b01100110; // b  **  **
			11'h13c: data_out = 8'b00000000; // c
			11'h13d: data_out = 8'b00000000; // d
			11'h13e: data_out = 8'b00000000; // e
			11'h13f: data_out = 8'b00000000; // f
			// code x14
			11'h140: data_out = 8'b00000000; // 0
			11'h141: data_out = 8'b00000000; // 1
			11'h142: data_out = 8'b01111111; // 2  *******
			11'h143: data_out = 8'b11011011; // 3 ** ** **
			11'h144: data_out = 8'b11011011; // 4 ** ** **
			11'h145: data_out = 8'b11011011; // 5 ** ** **
			11'h146: data_out = 8'b01111011; // 6  **** **
			11'h147: data_out = 8'b00011011; // 7    ** **
			11'h148: data_out = 8'b00011011; // 8    ** **
			11'h149: data_out = 8'b00011011; // 9    ** **
			11'h14a: data_out = 8'b00011011; // a    ** **
			11'h14b: data_out = 8'b00011011; // b    ** **
			11'h14c: data_out = 8'b00000000; // c
			11'h14d: data_out = 8'b00000000; // d
			11'h14e: data_out = 8'b00000000; // e
			11'h14f: data_out = 8'b00000000; // f
			// code x15
			11'h150: data_out = 8'b00000000; // 0
			11'h151: data_out = 8'b01111100; // 1  *****
			11'h152: data_out = 8'b11000110; // 2 **   **
			11'h153: data_out = 8'b01100000; // 3  **
			11'h154: data_out = 8'b00111000; // 4   ***
			11'h155: data_out = 8'b01101100; // 5  ** **
			11'h156: data_out = 8'b11000110; // 6 **   **
			11'h157: data_out = 8'b11000110; // 7 **   **
			11'h158: data_out = 8'b01101100; // 8  ** **
			11'h159: data_out = 8'b00111000; // 9   ***
			11'h15a: data_out = 8'b00001100; // a     **
			11'h15b: data_out = 8'b11000110; // b **   **
			11'h15c: data_out = 8'b01111100; // c  *****
			11'h15d: data_out = 8'b00000000; // d
			11'h15e: data_out = 8'b00000000; // e
			11'h15f: data_out = 8'b00000000; // f
			// code x16
			11'h160: data_out = 8'b00000000; // 0
			11'h161: data_out = 8'b00000000; // 1
			11'h162: data_out = 8'b00000000; // 2
			11'h163: data_out = 8'b00000000; // 3
			11'h164: data_out = 8'b00000000; // 4
			11'h165: data_out = 8'b00000000; // 5
			11'h166: data_out = 8'b00000000; // 6
			11'h167: data_out = 8'b00000000; // 7
			11'h168: data_out = 8'b11111110; // 8 *******
			11'h169: data_out = 8'b11111110; // 9 *******
			11'h16a: data_out = 8'b11111110; // a *******
			11'h16b: data_out = 8'b11111110; // b *******
			11'h16c: data_out = 8'b00000000; // c
			11'h16d: data_out = 8'b00000000; // d
			11'h16e: data_out = 8'b00000000; // e
			11'h16f: data_out = 8'b00000000; // f
			// code x17
			11'h170: data_out = 8'b00000000; // 0
			11'h171: data_out = 8'b00000000; // 1
			11'h172: data_out = 8'b00011000; // 2    **
			11'h173: data_out = 8'b00111100; // 3   ****
			11'h174: data_out = 8'b01111110; // 4  ******
			11'h175: data_out = 8'b00011000; // 5    **
			11'h176: data_out = 8'b00011000; // 6    **
			11'h177: data_out = 8'b00011000; // 7    **
			11'h178: data_out = 8'b01111110; // 8  ******
			11'h179: data_out = 8'b00111100; // 9   ****
			11'h17a: data_out = 8'b00011000; // a    **
			11'h17b: data_out = 8'b01111110; // b  ******
			11'h17c: data_out = 8'b00110000; // c
			11'h17d: data_out = 8'b00000000; // d
			11'h17e: data_out = 8'b00000000; // e
			11'h17f: data_out = 8'b00000000; // f
			// code x18
			11'h180: data_out = 8'b00000000; // 0
			11'h181: data_out = 8'b00000000; // 1
			11'h182: data_out = 8'b00011000; // 2    **
			11'h183: data_out = 8'b00111100; // 3   ****
			11'h184: data_out = 8'b01111110; // 4  ******
			11'h185: data_out = 8'b00011000; // 5    **
			11'h186: data_out = 8'b00011000; // 6    **
			11'h187: data_out = 8'b00011000; // 7    **
			11'h188: data_out = 8'b00011000; // 8    **
			11'h189: data_out = 8'b00011000; // 9    **
			11'h18a: data_out = 8'b00011000; // a    **
			11'h18b: data_out = 8'b00011000; // b    **
			11'h18c: data_out = 8'b00000000; // c
			11'h18d: data_out = 8'b00000000; // d
			11'h18e: data_out = 8'b00000000; // e
			11'h18f: data_out = 8'b00000000; // f
			// code x19
			11'h190: data_out = 8'b00000000; // 0
			11'h191: data_out = 8'b00000000; // 1
			11'h192: data_out = 8'b00011000; // 2    **
			11'h193: data_out = 8'b00011000; // 3    **
			11'h194: data_out = 8'b00011000; // 4    **
			11'h195: data_out = 8'b00011000; // 5    **
			11'h196: data_out = 8'b00011000; // 6    **
			11'h197: data_out = 8'b00011000; // 7    **
			11'h198: data_out = 8'b00011000; // 8    **
			11'h199: data_out = 8'b01111110; // 9  ******
			11'h19a: data_out = 8'b00111100; // a   ****
			11'h19b: data_out = 8'b00011000; // b    **
			11'h19c: data_out = 8'b00000000; // c
			11'h19d: data_out = 8'b00000000; // d
			11'h19e: data_out = 8'b00000000; // e
			11'h19f: data_out = 8'b00000000; // f
			// code x1a
			11'h1a0: data_out = 8'b00000000; // 0
			11'h1a1: data_out = 8'b00000000; // 1
			11'h1a2: data_out = 8'b00000000; // 2
			11'h1a3: data_out = 8'b00000000; // 3
			11'h1a4: data_out = 8'b00000000; // 4
			11'h1a5: data_out = 8'b00011000; // 5    **
			11'h1a6: data_out = 8'b00001100; // 6     **
			11'h1a7: data_out = 8'b11111110; // 7 *******
			11'h1a8: data_out = 8'b00001100; // 8     **
			11'h1a9: data_out = 8'b00011000; // 9    **
			11'h1aa: data_out = 8'b00000000; // a
			11'h1ab: data_out = 8'b00000000; // b
			11'h1ac: data_out = 8'b00000000; // c
			11'h1ad: data_out = 8'b00000000; // d
			11'h1ae: data_out = 8'b00000000; // e
			11'h1af: data_out = 8'b00000000; // f
			// code x1b
			11'h1b0: data_out = 8'b00000000; // 0
			11'h1b1: data_out = 8'b00000000; // 1
			11'h1b2: data_out = 8'b00000000; // 2
			11'h1b3: data_out = 8'b00000000; // 3
			11'h1b4: data_out = 8'b00000000; // 4
			11'h1b5: data_out = 8'b00110000; // 5   **
			11'h1b6: data_out = 8'b01100000; // 6  **
			11'h1b7: data_out = 8'b11111110; // 7 *******
			11'h1b8: data_out = 8'b01100000; // 8  **
			11'h1b9: data_out = 8'b00110000; // 9   **
			11'h1ba: data_out = 8'b00000000; // a
			11'h1bb: data_out = 8'b00000000; // b
			11'h1bc: data_out = 8'b00000000; // c
			11'h1bd: data_out = 8'b00000000; // d
			11'h1be: data_out = 8'b00000000; // e
			11'h1bf: data_out = 8'b00000000; // f
			// code x1c
			11'h1c0: data_out = 8'b00000000; // 0
			11'h1c1: data_out = 8'b00000000; // 1
			11'h1c2: data_out = 8'b00000000; // 2
			11'h1c3: data_out = 8'b00000000; // 3
			11'h1c4: data_out = 8'b00000000; // 4
			11'h1c5: data_out = 8'b00000000; // 5
			11'h1c6: data_out = 8'b11000000; // 6 **
			11'h1c7: data_out = 8'b11000000; // 7 **
			11'h1c8: data_out = 8'b11000000; // 8 **
			11'h1c9: data_out = 8'b11111110; // 9 *******
			11'h1ca: data_out = 8'b00000000; // a
			11'h1cb: data_out = 8'b00000000; // b
			11'h1cc: data_out = 8'b00000000; // c
			11'h1cd: data_out = 8'b00000000; // d
			11'h1ce: data_out = 8'b00000000; // e
			11'h1cf: data_out = 8'b00000000; // f
			// code x1d
			11'h1d0: data_out = 8'b00000000; // 0
			11'h1d1: data_out = 8'b00000000; // 1
			11'h1d2: data_out = 8'b00000000; // 2
			11'h1d3: data_out = 8'b00000000; // 3
			11'h1d4: data_out = 8'b00000000; // 4
			11'h1d5: data_out = 8'b00100100; // 5   *  *
			11'h1d6: data_out = 8'b01100110; // 6  **  **
			11'h1d7: data_out = 8'b11111111; // 7 ********
			11'h1d8: data_out = 8'b01100110; // 8  **  **
			11'h1d9: data_out = 8'b00100100; // 9   *  *
			11'h1da: data_out = 8'b00000000; // a
			11'h1db: data_out = 8'b00000000; // b
			11'h1dc: data_out = 8'b00000000; // c
			11'h1dd: data_out = 8'b00000000; // d
			11'h1de: data_out = 8'b00000000; // e
			11'h1df: data_out = 8'b00000000; // f
			// code x1e
			11'h1e0: data_out = 8'b00000000; // 0
			11'h1e1: data_out = 8'b00000000; // 1
			11'h1e2: data_out = 8'b00000000; // 2
			11'h1e3: data_out = 8'b00000000; // 3
			11'h1e4: data_out = 8'b00010000; // 4    *
			11'h1e5: data_out = 8'b00111000; // 5   ***
			11'h1e6: data_out = 8'b00111000; // 6   ***
			11'h1e7: data_out = 8'b01111100; // 7  *****
			11'h1e8: data_out = 8'b01111100; // 8  *****
			11'h1e9: data_out = 8'b11111110; // 9 *******
			11'h1ea: data_out = 8'b11111110; // a *******
			11'h1eb: data_out = 8'b00000000; // b
			11'h1ec: data_out = 8'b00000000; // c
			11'h1ed: data_out = 8'b00000000; // d
			11'h1ee: data_out = 8'b00000000; // e
			11'h1ef: data_out = 8'b00000000; // f
			// code x1f
			11'h1f0: data_out = 8'b00000000; // 0
			11'h1f1: data_out = 8'b00000000; // 1
			11'h1f2: data_out = 8'b00000000; // 2
			11'h1f3: data_out = 8'b00000000; // 3
			11'h1f4: data_out = 8'b11111110; // 4 *******
			11'h1f5: data_out = 8'b11111110; // 5 *******
			11'h1f6: data_out = 8'b01111100; // 6  *****
			11'h1f7: data_out = 8'b01111100; // 7  *****
			11'h1f8: data_out = 8'b00111000; // 8   ***
			11'h1f9: data_out = 8'b00111000; // 9   ***
			11'h1fa: data_out = 8'b00010000; // a    *
			11'h1fb: data_out = 8'b00000000; // b
			11'h1fc: data_out = 8'b00000000; // c
			11'h1fd: data_out = 8'b00000000; // d
			11'h1fe: data_out = 8'b00000000; // e
			11'h1ff: data_out = 8'b00000000; // f
			// code x20
			11'h200: data_out = 8'b00000000; // 0
			11'h201: data_out = 8'b00000000; // 1
			11'h202: data_out = 8'b00000000; // 2
			11'h203: data_out = 8'b00000000; // 3
			11'h204: data_out = 8'b00000000; // 4
			11'h205: data_out = 8'b00000000; // 5
			11'h206: data_out = 8'b00000000; // 6
			11'h207: data_out = 8'b00000000; // 7
			11'h208: data_out = 8'b00000000; // 8
			11'h209: data_out = 8'b00000000; // 9
			11'h20a: data_out = 8'b00000000; // a
			11'h20b: data_out = 8'b00000000; // b
			11'h20c: data_out = 8'b00000000; // c
			11'h20d: data_out = 8'b00000000; // d
			11'h20e: data_out = 8'b00000000; // e
			11'h20f: data_out = 8'b00000000; // f
			// code x21
			11'h210: data_out = 8'b00000000; // 0
			11'h211: data_out = 8'b00000000; // 1
			11'h212: data_out = 8'b00011000; // 2    **
			11'h213: data_out = 8'b00111100; // 3   ****
			11'h214: data_out = 8'b00111100; // 4   ****
			11'h215: data_out = 8'b00111100; // 5   ****
			11'h216: data_out = 8'b00011000; // 6    **
			11'h217: data_out = 8'b00011000; // 7    **
			11'h218: data_out = 8'b00011000; // 8    **
			11'h219: data_out = 8'b00000000; // 9
			11'h21a: data_out = 8'b00011000; // a    **
			11'h21b: data_out = 8'b00011000; // b    **
			11'h21c: data_out = 8'b00000000; // c
			11'h21d: data_out = 8'b00000000; // d
			11'h21e: data_out = 8'b00000000; // e
			11'h21f: data_out = 8'b00000000; // f
			// code x22
			11'h220: data_out = 8'b00000000; // 0
			11'h221: data_out = 8'b01100110; // 1  **  **
			11'h222: data_out = 8'b01100110; // 2  **  **
			11'h223: data_out = 8'b01100110; // 3  **  **
			11'h224: data_out = 8'b00100100; // 4   *  *
			11'h225: data_out = 8'b00000000; // 5
			11'h226: data_out = 8'b00000000; // 6
			11'h227: data_out = 8'b00000000; // 7
			11'h228: data_out = 8'b00000000; // 8
			11'h229: data_out = 8'b00000000; // 9
			11'h22a: data_out = 8'b00000000; // a
			11'h22b: data_out = 8'b00000000; // b
			11'h22c: data_out = 8'b00000000; // c
			11'h22d: data_out = 8'b00000000; // d
			11'h22e: data_out = 8'b00000000; // e
			11'h22f: data_out = 8'b00000000; // f
			// code x23
			11'h230: data_out = 8'b00000000; // 0
			11'h231: data_out = 8'b00000000; // 1
			11'h232: data_out = 8'b00000000; // 2
			11'h233: data_out = 8'b01101100; // 3  ** **
			11'h234: data_out = 8'b01101100; // 4  ** **
			11'h235: data_out = 8'b11111110; // 5 *******
			11'h236: data_out = 8'b01101100; // 6  ** **
			11'h237: data_out = 8'b01101100; // 7  ** **
			11'h238: data_out = 8'b01101100; // 8  ** **
			11'h239: data_out = 8'b11111110; // 9 *******
			11'h23a: data_out = 8'b01101100; // a  ** **
			11'h23b: data_out = 8'b01101100; // b  ** **
			11'h23c: data_out = 8'b00000000; // c
			11'h23d: data_out = 8'b00000000; // d
			11'h23e: data_out = 8'b00000000; // e
			11'h23f: data_out = 8'b00000000; // f
			// code x24
			11'h240: data_out = 8'b00011000; // 0     **
			11'h241: data_out = 8'b00011000; // 1     **
			11'h242: data_out = 8'b01111100; // 2   *****
			11'h243: data_out = 8'b11000110; // 3  **   **
			11'h244: data_out = 8'b11000010; // 4  **    *
			11'h245: data_out = 8'b11000000; // 5  **
			11'h246: data_out = 8'b01111100; // 6   *****
			11'h247: data_out = 8'b00000110; // 7       **
			11'h248: data_out = 8'b00000110; // 8       **
			11'h249: data_out = 8'b10000110; // 9  *    **
			11'h24a: data_out = 8'b11000110; // a  **   **
			11'h24b: data_out = 8'b01111100; // b   *****
			11'h24c: data_out = 8'b00011000; // c     **
			11'h24d: data_out = 8'b00011000; // d     **
			11'h24e: data_out = 8'b00000000; // e
			11'h24f: data_out = 8'b00000000; // f
			// code x25
			11'h250: data_out = 8'b00000000; // 0
			11'h251: data_out = 8'b00000000; // 1
			11'h252: data_out = 8'b00000000; // 2
			11'h253: data_out = 8'b00000000; // 3
			11'h254: data_out = 8'b11000010; // 4 **    *
			11'h255: data_out = 8'b11000110; // 5 **   **
			11'h256: data_out = 8'b00001100; // 6     **
			11'h257: data_out = 8'b00011000; // 7    **
			11'h258: data_out = 8'b00110000; // 8   **
			11'h259: data_out = 8'b01100000; // 9  **
			11'h25a: data_out = 8'b11000110; // a **   **
			11'h25b: data_out = 8'b10000110; // b *    **
			11'h25c: data_out = 8'b00000000; // c
			11'h25d: data_out = 8'b00000000; // d
			11'h25e: data_out = 8'b00000000; // e
			11'h25f: data_out = 8'b00000000; // f
			// code x26
			11'h260: data_out = 8'b00000000; // 0
			11'h261: data_out = 8'b00000000; // 1
			11'h262: data_out = 8'b00111000; // 2   ***
			11'h263: data_out = 8'b01101100; // 3  ** **
			11'h264: data_out = 8'b01101100; // 4  ** **
			11'h265: data_out = 8'b00111000; // 5   ***
			11'h266: data_out = 8'b01110110; // 6  *** **
			11'h267: data_out = 8'b11011100; // 7 ** ***
			11'h268: data_out = 8'b11001100; // 8 **  **
			11'h269: data_out = 8'b11001100; // 9 **  **
			11'h26a: data_out = 8'b11001100; // a **  **
			11'h26b: data_out = 8'b01110110; // b  *** **
			11'h26c: data_out = 8'b00000000; // c
			11'h26d: data_out = 8'b00000000; // d
			11'h26e: data_out = 8'b00000000; // e
			11'h26f: data_out = 8'b00000000; // f
			// code x27
			11'h270: data_out = 8'b00000000; // 0
			11'h271: data_out = 8'b00110000; // 1   **
			11'h272: data_out = 8'b00110000; // 2   **
			11'h273: data_out = 8'b00110000; // 3   **
			11'h274: data_out = 8'b01100000; // 4  **
			11'h275: data_out = 8'b00000000; // 5
			11'h276: data_out = 8'b00000000; // 6
			11'h277: data_out = 8'b00000000; // 7
			11'h278: data_out = 8'b00000000; // 8
			11'h279: data_out = 8'b00000000; // 9
			11'h27a: data_out = 8'b00000000; // a
			11'h27b: data_out = 8'b00000000; // b
			11'h27c: data_out = 8'b00000000; // c
			11'h27d: data_out = 8'b00000000; // d
			11'h27e: data_out = 8'b00000000; // e
			11'h27f: data_out = 8'b00000000; // f
			// code x28
			11'h280: data_out = 8'b00000000; // 0
			11'h281: data_out = 8'b00000000; // 1
			11'h282: data_out = 8'b00001100; // 2     **
			11'h283: data_out = 8'b00011000; // 3    **
			11'h284: data_out = 8'b00110000; // 4   **
			11'h285: data_out = 8'b00110000; // 5   **
			11'h286: data_out = 8'b00110000; // 6   **
			11'h287: data_out = 8'b00110000; // 7   **
			11'h288: data_out = 8'b00110000; // 8   **
			11'h289: data_out = 8'b00110000; // 9   **
			11'h28a: data_out = 8'b00011000; // a    **
			11'h28b: data_out = 8'b00001100; // b     **
			11'h28c: data_out = 8'b00000000; // c
			11'h28d: data_out = 8'b00000000; // d
			11'h28e: data_out = 8'b00000000; // e
			11'h28f: data_out = 8'b00000000; // f
			// code x29
			11'h290: data_out = 8'b00000000; // 0
			11'h291: data_out = 8'b00000000; // 1
			11'h292: data_out = 8'b00110000; // 2   **
			11'h293: data_out = 8'b00011000; // 3    **
			11'h294: data_out = 8'b00001100; // 4     **
			11'h295: data_out = 8'b00001100; // 5     **
			11'h296: data_out = 8'b00001100; // 6     **
			11'h297: data_out = 8'b00001100; // 7     **
			11'h298: data_out = 8'b00001100; // 8     **
			11'h299: data_out = 8'b00001100; // 9     **
			11'h29a: data_out = 8'b00011000; // a    **
			11'h29b: data_out = 8'b00110000; // b   **
			11'h29c: data_out = 8'b00000000; // c
			11'h29d: data_out = 8'b00000000; // d
			11'h29e: data_out = 8'b00000000; // e
			11'h29f: data_out = 8'b00000000; // f
			// code x2a
			11'h2a0: data_out = 8'b00000000; // 0
			11'h2a1: data_out = 8'b00000000; // 1
			11'h2a2: data_out = 8'b00000000; // 2
			11'h2a3: data_out = 8'b00000000; // 3
			11'h2a4: data_out = 8'b00000000; // 4
			11'h2a5: data_out = 8'b01100110; // 5  **  **
			11'h2a6: data_out = 8'b00111100; // 6   ****
			11'h2a7: data_out = 8'b11111111; // 7 ********
			11'h2a8: data_out = 8'b00111100; // 8   ****
			11'h2a9: data_out = 8'b01100110; // 9  **  **
			11'h2aa: data_out = 8'b00000000; // a
			11'h2ab: data_out = 8'b00000000; // b
			11'h2ac: data_out = 8'b00000000; // c
			11'h2ad: data_out = 8'b00000000; // d
			11'h2ae: data_out = 8'b00000000; // e
			11'h2af: data_out = 8'b00000000; // f
			// code x2b
			11'h2b0: data_out = 8'b00000000; // 0
			11'h2b1: data_out = 8'b00000000; // 1
			11'h2b2: data_out = 8'b00000000; // 2
			11'h2b3: data_out = 8'b00000000; // 3
			11'h2b4: data_out = 8'b00000000; // 4
			11'h2b5: data_out = 8'b00011000; // 5    **
			11'h2b6: data_out = 8'b00011000; // 6    **
			11'h2b7: data_out = 8'b01111110; // 7  ******
			11'h2b8: data_out = 8'b00011000; // 8    **
			11'h2b9: data_out = 8'b00011000; // 9    **
			11'h2ba: data_out = 8'b00000000; // a
			11'h2bb: data_out = 8'b00000000; // b
			11'h2bc: data_out = 8'b00000000; // c
			11'h2bd: data_out = 8'b00000000; // d
			11'h2be: data_out = 8'b00000000; // e
			11'h2bf: data_out = 8'b00000000; // f
			// code x2c
			11'h2c0: data_out = 8'b00000000; // 0
			11'h2c1: data_out = 8'b00000000; // 1
			11'h2c2: data_out = 8'b00000000; // 2
			11'h2c3: data_out = 8'b00000000; // 3
			11'h2c4: data_out = 8'b00000000; // 4
			11'h2c5: data_out = 8'b00000000; // 5
			11'h2c6: data_out = 8'b00000000; // 6
			11'h2c7: data_out = 8'b00000000; // 7
			11'h2c8: data_out = 8'b00000000; // 8
			11'h2c9: data_out = 8'b00011000; // 9    **
			11'h2ca: data_out = 8'b00011000; // a    **
			11'h2cb: data_out = 8'b00011000; // b    **
			11'h2cc: data_out = 8'b00110000; // c   **
			11'h2cd: data_out = 8'b00000000; // d
			11'h2ce: data_out = 8'b00000000; // e
			11'h2cf: data_out = 8'b00000000; // f
			// code x2d
			11'h2d0: data_out = 8'b00000000; // 0
			11'h2d1: data_out = 8'b00000000; // 1
			11'h2d2: data_out = 8'b00000000; // 2
			11'h2d3: data_out = 8'b00000000; // 3
			11'h2d4: data_out = 8'b00000000; // 4
			11'h2d5: data_out = 8'b00000000; // 5
			11'h2d6: data_out = 8'b00000000; // 6
			11'h2d7: data_out = 8'b01111110; // 7  ******
			11'h2d8: data_out = 8'b00000000; // 8
			11'h2d9: data_out = 8'b00000000; // 9
			11'h2da: data_out = 8'b00000000; // a
			11'h2db: data_out = 8'b00000000; // b
			11'h2dc: data_out = 8'b00000000; // c
			11'h2dd: data_out = 8'b00000000; // d
			11'h2de: data_out = 8'b00000000; // e
			11'h2df: data_out = 8'b00000000; // f
			// code x2e
			11'h2e0: data_out = 8'b00000000; // 0
			11'h2e1: data_out = 8'b00000000; // 1
			11'h2e2: data_out = 8'b00000000; // 2
			11'h2e3: data_out = 8'b00000000; // 3
			11'h2e4: data_out = 8'b00000000; // 4
			11'h2e5: data_out = 8'b00000000; // 5
			11'h2e6: data_out = 8'b00000000; // 6
			11'h2e7: data_out = 8'b00000000; // 7
			11'h2e8: data_out = 8'b00000000; // 8
			11'h2e9: data_out = 8'b00000000; // 9
			11'h2ea: data_out = 8'b00011000; // a    **
			11'h2eb: data_out = 8'b00011000; // b    **
			11'h2ec: data_out = 8'b00000000; // c
			11'h2ed: data_out = 8'b00000000; // d
			11'h2ee: data_out = 8'b00000000; // e
			11'h2ef: data_out = 8'b00000000; // f
			// code x2f
			11'h2f0: data_out = 8'b00000000; // 0
			11'h2f1: data_out = 8'b00000000; // 1
			11'h2f2: data_out = 8'b00000000; // 2
			11'h2f3: data_out = 8'b00000000; // 3
			11'h2f4: data_out = 8'b00000010; // 4       *
			11'h2f5: data_out = 8'b00000110; // 5      **
			11'h2f6: data_out = 8'b00001100; // 6     **
			11'h2f7: data_out = 8'b00011000; // 7    **
			11'h2f8: data_out = 8'b00110000; // 8   **
			11'h2f9: data_out = 8'b01100000; // 9  **
			11'h2fa: data_out = 8'b11000000; // a **
			11'h2fb: data_out = 8'b10000000; // b *
			11'h2fc: data_out = 8'b00000000; // c
			11'h2fd: data_out = 8'b00000000; // d
			11'h2fe: data_out = 8'b00000000; // e
			11'h2ff: data_out = 8'b00000000; // f
			// code x30
			11'h300: data_out = 8'b00000000; // 0
			11'h301: data_out = 8'b00000000; // 1
			11'h302: data_out = 8'b01111100; // 2  *****
			11'h303: data_out = 8'b11000110; // 3 **   **
			11'h304: data_out = 8'b11000110; // 4 **   **
			11'h305: data_out = 8'b11001110; // 5 **  ***
			11'h306: data_out = 8'b11011110; // 6 ** ****
			11'h307: data_out = 8'b11110110; // 7 **** **
			11'h308: data_out = 8'b11100110; // 8 ***  **
			11'h309: data_out = 8'b11000110; // 9 **   **
			11'h30a: data_out = 8'b11000110; // a **   **
			11'h30b: data_out = 8'b01111100; // b  *****
			11'h30c: data_out = 8'b00000000; // c
			11'h30d: data_out = 8'b00000000; // d
			11'h30e: data_out = 8'b00000000; // e
			11'h30f: data_out = 8'b00000000; // f
			// code x31
			11'h310: data_out = 8'b00000000; // 0
			11'h311: data_out = 8'b00000000; // 1
			11'h312: data_out = 8'b00011000; // 2    **
			11'h313: data_out = 8'b00111000; // 3   ***
			11'h314: data_out = 8'b01111000; // 4  ****
			11'h315: data_out = 8'b00011000; // 5    **
			11'h316: data_out = 8'b00011000; // 6    **
			11'h317: data_out = 8'b00011000; // 7    **
			11'h318: data_out = 8'b00011000; // 8    **
			11'h319: data_out = 8'b00011000; // 9    **
			11'h31a: data_out = 8'b00011000; // a    **
			11'h31b: data_out = 8'b01111110; // b  ******
			11'h31c: data_out = 8'b00000000; // c    
			11'h31d: data_out = 8'b00000000; // d
			11'h31e: data_out = 8'b00000000; // e
			11'h31f: data_out = 8'b00000000; // f
			// code x32
			11'h320: data_out = 8'b00000000; // 0
			11'h321: data_out = 8'b00000000; // 1
			11'h322: data_out = 8'b01111100; // 2  *****
			11'h323: data_out = 8'b11000110; // 3 **   **
			11'h324: data_out = 8'b00000110; // 4      **
			11'h325: data_out = 8'b00001100; // 5     **
			11'h326: data_out = 8'b00011000; // 6    **
			11'h327: data_out = 8'b00110000; // 7   **
			11'h328: data_out = 8'b01100000; // 8  **
			11'h329: data_out = 8'b11000000; // 9 **
			11'h32a: data_out = 8'b11000110; // a **   **
			11'h32b: data_out = 8'b11111110; // b *******
			11'h32c: data_out = 8'b00000000; // c
			11'h32d: data_out = 8'b00000000; // d
			11'h32e: data_out = 8'b00000000; // e
			11'h32f: data_out = 8'b00000000; // f
			// code x33
			11'h330: data_out = 8'b00000000; // 0
			11'h331: data_out = 8'b00000000; // 1
			11'h332: data_out = 8'b01111100; // 2  *****
			11'h333: data_out = 8'b11000110; // 3 **   **
			11'h334: data_out = 8'b00000110; // 4      **
			11'h335: data_out = 8'b00000110; // 5      **
			11'h336: data_out = 8'b00111100; // 6   ****
			11'h337: data_out = 8'b00000110; // 7      **
			11'h338: data_out = 8'b00000110; // 8      **
			11'h339: data_out = 8'b00000110; // 9      **
			11'h33a: data_out = 8'b11000110; // a **   **
			11'h33b: data_out = 8'b01111100; // b  *****
			11'h33c: data_out = 8'b00000000; // c
			11'h33d: data_out = 8'b00000000; // d
			11'h33e: data_out = 8'b00000000; // e
			11'h33f: data_out = 8'b00000000; // f
			// code x34
			11'h340: data_out = 8'b00000000; // 0
			11'h341: data_out = 8'b00000000; // 1
			11'h342: data_out = 8'b00001100; // 2     **
			11'h343: data_out = 8'b00011100; // 3    ***
			11'h344: data_out = 8'b00111100; // 4   ****
			11'h345: data_out = 8'b01101100; // 5  ** **
			11'h346: data_out = 8'b11001100; // 6 **  **
			11'h347: data_out = 8'b11111110; // 7 *******
			11'h348: data_out = 8'b00001100; // 8     **
			11'h349: data_out = 8'b00001100; // 9     **
			11'h34a: data_out = 8'b00001100; // a     **
			11'h34b: data_out = 8'b00011110; // b    ****
			11'h34c: data_out = 8'b00000000; // c
			11'h34d: data_out = 8'b00000000; // d
			11'h34e: data_out = 8'b00000000; // e
			11'h34f: data_out = 8'b00000000; // f
			// code x35
			11'h350: data_out = 8'b00000000; // 0
			11'h351: data_out = 8'b00000000; // 1
			11'h352: data_out = 8'b11111110; // 2 *******
			11'h353: data_out = 8'b11000000; // 3 **
			11'h354: data_out = 8'b11000000; // 4 **
			11'h355: data_out = 8'b11000000; // 5 **
			11'h356: data_out = 8'b11111100; // 6 ******
			11'h357: data_out = 8'b00000110; // 7      **
			11'h358: data_out = 8'b00000110; // 8      **
			11'h359: data_out = 8'b00000110; // 9      **
			11'h35a: data_out = 8'b11000110; // a **   **
			11'h35b: data_out = 8'b01111100; // b  *****
			11'h35c: data_out = 8'b00000000; // c
			11'h35d: data_out = 8'b00000000; // d
			11'h35e: data_out = 8'b00000000; // e
			11'h35f: data_out = 8'b00000000; // f
			// code x36
			11'h360: data_out = 8'b00000000; // 0
			11'h361: data_out = 8'b00000000; // 1
			11'h362: data_out = 8'b00111000; // 2   ***
			11'h363: data_out = 8'b01100000; // 3  **
			11'h364: data_out = 8'b11000000; // 4 **
			11'h365: data_out = 8'b11000000; // 5 **
			11'h366: data_out = 8'b11111100; // 6 ******
			11'h367: data_out = 8'b11000110; // 7 **   **
			11'h368: data_out = 8'b11000110; // 8 **   **
			11'h369: data_out = 8'b11000110; // 9 **   **
			11'h36a: data_out = 8'b11000110; // a **   **
			11'h36b: data_out = 8'b01111100; // b  *****
			11'h36c: data_out = 8'b00000000; // c
			11'h36d: data_out = 8'b00000000; // d
			11'h36e: data_out = 8'b00000000; // e
			11'h36f: data_out = 8'b00000000; // f
			// code x37
			11'h370: data_out = 8'b00000000; // 0
			11'h371: data_out = 8'b00000000; // 1
			11'h372: data_out = 8'b11111110; // 2 *******
			11'h373: data_out = 8'b11000110; // 3 **   **
			11'h374: data_out = 8'b00000110; // 4      **
			11'h375: data_out = 8'b00000110; // 5      **
			11'h376: data_out = 8'b00001100; // 6     **
			11'h377: data_out = 8'b00011000; // 7    **
			11'h378: data_out = 8'b00110000; // 8   **
			11'h379: data_out = 8'b00110000; // 9   **
			11'h37a: data_out = 8'b00110000; // a   **
			11'h37b: data_out = 8'b00110000; // b   **
			11'h37c: data_out = 8'b00000000; // c
			11'h37d: data_out = 8'b00000000; // d
			11'h37e: data_out = 8'b00000000; // e
			11'h37f: data_out = 8'b00000000; // f
			// code x38
			11'h380: data_out = 8'b00000000; // 0
			11'h381: data_out = 8'b00000000; // 1
			11'h382: data_out = 8'b01111100; // 2  *****
			11'h383: data_out = 8'b11000110; // 3 **   **
			11'h384: data_out = 8'b11000110; // 4 **   **
			11'h385: data_out = 8'b11000110; // 5 **   **
			11'h386: data_out = 8'b01111100; // 6  *****
			11'h387: data_out = 8'b11000110; // 7 **   **
			11'h388: data_out = 8'b11000110; // 8 **   **
			11'h389: data_out = 8'b11000110; // 9 **   **
			11'h38a: data_out = 8'b11000110; // a **   **
			11'h38b: data_out = 8'b01111100; // b  *****
			11'h38c: data_out = 8'b00000000; // c
			11'h38d: data_out = 8'b00000000; // d
			11'h38e: data_out = 8'b00000000; // e
			11'h38f: data_out = 8'b00000000; // f
			// code x39
			11'h390: data_out = 8'b00000000; // 0
			11'h391: data_out = 8'b00000000; // 1
			11'h392: data_out = 8'b01111100; // 2  *****
			11'h393: data_out = 8'b11000110; // 3 **   **
			11'h394: data_out = 8'b11000110; // 4 **   **
			11'h395: data_out = 8'b11000110; // 5 **   **
			11'h396: data_out = 8'b01111110; // 6  ******
			11'h397: data_out = 8'b00000110; // 7      **
			11'h398: data_out = 8'b00000110; // 8      **
			11'h399: data_out = 8'b00000110; // 9      **
			11'h39a: data_out = 8'b00001100; // a     **
			11'h39b: data_out = 8'b01111000; // b  ****
			11'h39c: data_out = 8'b00000000; // c
			11'h39d: data_out = 8'b00000000; // d
			11'h39e: data_out = 8'b00000000; // e
			11'h39f: data_out = 8'b00000000; // f
			// code x3a
			11'h3a0: data_out = 8'b00000000; // 0
			11'h3a1: data_out = 8'b00000000; // 1
			11'h3a2: data_out = 8'b00000000; // 2
			11'h3a3: data_out = 8'b00000000; // 3
			11'h3a4: data_out = 8'b00011000; // 4    **
			11'h3a5: data_out = 8'b00011000; // 5    **
			11'h3a6: data_out = 8'b00000000; // 6
			11'h3a7: data_out = 8'b00000000; // 7
			11'h3a8: data_out = 8'b00000000; // 8
			11'h3a9: data_out = 8'b00011000; // 9    **
			11'h3aa: data_out = 8'b00011000; // a    **
			11'h3ab: data_out = 8'b00000000; // b
			11'h3ac: data_out = 8'b00000000; // c
			11'h3ad: data_out = 8'b00000000; // d
			11'h3ae: data_out = 8'b00000000; // e
			11'h3af: data_out = 8'b00000000; // f
			// code x3b
			11'h3b0: data_out = 8'b00000000; // 0
			11'h3b1: data_out = 8'b00000000; // 1
			11'h3b2: data_out = 8'b00000000; // 2
			11'h3b3: data_out = 8'b00000000; // 3
			11'h3b4: data_out = 8'b00011000; // 4    **
			11'h3b5: data_out = 8'b00011000; // 5    **
			11'h3b6: data_out = 8'b00000000; // 6
			11'h3b7: data_out = 8'b00000000; // 7
			11'h3b8: data_out = 8'b00000000; // 8
			11'h3b9: data_out = 8'b00011000; // 9    **
			11'h3ba: data_out = 8'b00011000; // a    **
			11'h3bb: data_out = 8'b00110000; // b   **
			11'h3bc: data_out = 8'b00000000; // c
			11'h3bd: data_out = 8'b00000000; // d
			11'h3be: data_out = 8'b00000000; // e
			11'h3bf: data_out = 8'b00000000; // f
			// code x3c
			11'h3c0: data_out = 8'b00000000; // 0
			11'h3c1: data_out = 8'b00000000; // 1
			11'h3c2: data_out = 8'b00000000; // 2
			11'h3c3: data_out = 8'b00000110; // 3      **
			11'h3c4: data_out = 8'b00001100; // 4     **
			11'h3c5: data_out = 8'b00011000; // 5    **
			11'h3c6: data_out = 8'b00110000; // 6   **
			11'h3c7: data_out = 8'b01100000; // 7  **
			11'h3c8: data_out = 8'b00110000; // 8   **
			11'h3c9: data_out = 8'b00011000; // 9    **
			11'h3ca: data_out = 8'b00001100; // a     **
			11'h3cb: data_out = 8'b00000110; // b      **
			11'h3cc: data_out = 8'b00000000; // c
			11'h3cd: data_out = 8'b00000000; // d
			11'h3ce: data_out = 8'b00000000; // e
			11'h3cf: data_out = 8'b00000000; // f
			// code x3d
			11'h3d0: data_out = 8'b00000000; // 0
			11'h3d1: data_out = 8'b00000000; // 1
			11'h3d2: data_out = 8'b00000000; // 2
			11'h3d3: data_out = 8'b00000000; // 3
			11'h3d4: data_out = 8'b00000000; // 4
			11'h3d5: data_out = 8'b01111110; // 5  ******
			11'h3d6: data_out = 8'b00000000; // 6
			11'h3d7: data_out = 8'b00000000; // 7
			11'h3d8: data_out = 8'b01111110; // 8  ******
			11'h3d9: data_out = 8'b00000000; // 9
			11'h3da: data_out = 8'b00000000; // a
			11'h3db: data_out = 8'b00000000; // b
			11'h3dc: data_out = 8'b00000000; // c
			11'h3dd: data_out = 8'b00000000; // d
			11'h3de: data_out = 8'b00000000; // e
			11'h3df: data_out = 8'b00000000; // f
			// code x3e
			11'h3e0: data_out = 8'b00000000; // 0
			11'h3e1: data_out = 8'b00000000; // 1
			11'h3e2: data_out = 8'b00000000; // 2
			11'h3e3: data_out = 8'b01100000; // 3  **
			11'h3e4: data_out = 8'b00110000; // 4   **
			11'h3e5: data_out = 8'b00011000; // 5    **
			11'h3e6: data_out = 8'b00001100; // 6     **
			11'h3e7: data_out = 8'b00000110; // 7      **
			11'h3e8: data_out = 8'b00001100; // 8     **
			11'h3e9: data_out = 8'b00011000; // 9    **
			11'h3ea: data_out = 8'b00110000; // a   **
			11'h3eb: data_out = 8'b01100000; // b  **
			11'h3ec: data_out = 8'b00000000; // c
			11'h3ed: data_out = 8'b00000000; // d
			11'h3ee: data_out = 8'b00000000; // e
			11'h3ef: data_out = 8'b00000000; // f
			// code x3f
			11'h3f0: data_out = 8'b00000000; // 0
			11'h3f1: data_out = 8'b00000000; // 1
			11'h3f2: data_out = 8'b01111100; // 2  *****
			11'h3f3: data_out = 8'b11000110; // 3 **   **
			11'h3f4: data_out = 8'b11000110; // 4 **   **
			11'h3f5: data_out = 8'b00001100; // 5     **
			11'h3f6: data_out = 8'b00011000; // 6    **
			11'h3f7: data_out = 8'b00011000; // 7    **
			11'h3f8: data_out = 8'b00011000; // 8    **
			11'h3f9: data_out = 8'b00000000; // 9
			11'h3fa: data_out = 8'b00011000; // a    **
			11'h3fb: data_out = 8'b00011000; // b    **
			11'h3fc: data_out = 8'b00000000; // c
			11'h3fd: data_out = 8'b00000000; // d
			11'h3fe: data_out = 8'b00000000; // e
			11'h3ff: data_out = 8'b00000000; // f
			// code x40
			11'h400: data_out = 8'b00000000; // 0
			11'h401: data_out = 8'b00000000; // 1
			11'h402: data_out = 8'b01111100; // 2  *****
			11'h403: data_out = 8'b11000110; // 3 **   **
			11'h404: data_out = 8'b11000110; // 4 **   **
			11'h405: data_out = 8'b11000110; // 5 **   **
			11'h406: data_out = 8'b11011110; // 6 ** ****
			11'h407: data_out = 8'b11011110; // 7 ** ****
			11'h408: data_out = 8'b11011110; // 8 ** ****
			11'h409: data_out = 8'b11011100; // 9 ** ***
			11'h40a: data_out = 8'b11000000; // a **
			11'h40b: data_out = 8'b01111100; // b  *****
			11'h40c: data_out = 8'b00000000; // c
			11'h40d: data_out = 8'b00000000; // d
			11'h40e: data_out = 8'b00000000; // e
			11'h40f: data_out = 8'b00000000; // f
			// code x41
			11'h410: data_out = 8'b00000000; // 0
			11'h411: data_out = 8'b00000000; // 1
			11'h412: data_out = 8'b00010000; // 2    *
			11'h413: data_out = 8'b00111000; // 3   ***
			11'h414: data_out = 8'b01101100; // 4  ** **
			11'h415: data_out = 8'b11000110; // 5 **   **
			11'h416: data_out = 8'b11000110; // 6 **   **
			11'h417: data_out = 8'b11111110; // 7 *******
			11'h418: data_out = 8'b11000110; // 8 **   **
			11'h419: data_out = 8'b11000110; // 9 **   **
			11'h41a: data_out = 8'b11000110; // a **   **
			11'h41b: data_out = 8'b11000110; // b **   **
			11'h41c: data_out = 8'b00000000; // c
			11'h41d: data_out = 8'b00000000; // d
			11'h41e: data_out = 8'b00000000; // e
			11'h41f: data_out = 8'b00000000; // f
			// code x42
			11'h420: data_out = 8'b00000000; // 0
			11'h421: data_out = 8'b00000000; // 1
			11'h422: data_out = 8'b11111100; // 2 ******
			11'h423: data_out = 8'b01100110; // 3  **  **
			11'h424: data_out = 8'b01100110; // 4  **  **
			11'h425: data_out = 8'b01100110; // 5  **  **
			11'h426: data_out = 8'b01111100; // 6  *****
			11'h427: data_out = 8'b01100110; // 7  **  **
			11'h428: data_out = 8'b01100110; // 8  **  **
			11'h429: data_out = 8'b01100110; // 9  **  **
			11'h42a: data_out = 8'b01100110; // a  **  **
			11'h42b: data_out = 8'b11111100; // b ******
			11'h42c: data_out = 8'b00000000; // c
			11'h42d: data_out = 8'b00000000; // d
			11'h42e: data_out = 8'b00000000; // e
			11'h42f: data_out = 8'b00000000; // f
			// code x43
			11'h430: data_out = 8'b00000000; // 0
			11'h431: data_out = 8'b00000000; // 1
			11'h432: data_out = 8'b00111100; // 2   ****
			11'h433: data_out = 8'b01100110; // 3  **  **
			11'h434: data_out = 8'b11000010; // 4 **    *
			11'h435: data_out = 8'b11000000; // 5 **
			11'h436: data_out = 8'b11000000; // 6 **
			11'h437: data_out = 8'b11000000; // 7 **
			11'h438: data_out = 8'b11000000; // 8 **
			11'h439: data_out = 8'b11000010; // 9 **    *
			11'h43a: data_out = 8'b01100110; // a  **  **
			11'h43b: data_out = 8'b00111100; // b   ****
			11'h43c: data_out = 8'b00000000; // c
			11'h43d: data_out = 8'b00000000; // d
			11'h43e: data_out = 8'b00000000; // e
			11'h43f: data_out = 8'b00000000; // f
			// code x44
			11'h440: data_out = 8'b00000000; // 0
			11'h441: data_out = 8'b00000000; // 1
			11'h442: data_out = 8'b11111000; // 2 *****
			11'h443: data_out = 8'b01101100; // 3  ** **
			11'h444: data_out = 8'b01100110; // 4  **  **
			11'h445: data_out = 8'b01100110; // 5  **  **
			11'h446: data_out = 8'b01100110; // 6  **  **
			11'h447: data_out = 8'b01100110; // 7  **  **
			11'h448: data_out = 8'b01100110; // 8  **  **
			11'h449: data_out = 8'b01100110; // 9  **  **
			11'h44a: data_out = 8'b01101100; // a  ** **
			11'h44b: data_out = 8'b11111000; // b *****
			11'h44c: data_out = 8'b00000000; // c
			11'h44d: data_out = 8'b00000000; // d
			11'h44e: data_out = 8'b00000000; // e
			11'h44f: data_out = 8'b00000000; // f
			// code x45
			11'h450: data_out = 8'b00000000; // 0
			11'h451: data_out = 8'b00000000; // 1
			11'h452: data_out = 8'b11111110; // 2 *******
			11'h453: data_out = 8'b01100110; // 3  **  **
			11'h454: data_out = 8'b01100010; // 4  **   *
			11'h455: data_out = 8'b01101000; // 5  ** *
			11'h456: data_out = 8'b01111000; // 6  ****
			11'h457: data_out = 8'b01101000; // 7  ** *
			11'h458: data_out = 8'b01100000; // 8  **
			11'h459: data_out = 8'b01100010; // 9  **   *
			11'h45a: data_out = 8'b01100110; // a  **  **
			11'h45b: data_out = 8'b11111110; // b *******
			11'h45c: data_out = 8'b00000000; // c
			11'h45d: data_out = 8'b00000000; // d
			11'h45e: data_out = 8'b00000000; // e
			11'h45f: data_out = 8'b00000000; // f
			// code x46
			11'h460: data_out = 8'b00000000; // 0
			11'h461: data_out = 8'b00000000; // 1
			11'h462: data_out = 8'b11111110; // 2 *******
			11'h463: data_out = 8'b01100110; // 3  **  **
			11'h464: data_out = 8'b01100010; // 4  **   *
			11'h465: data_out = 8'b01101000; // 5  ** *
			11'h466: data_out = 8'b01111000; // 6  ****
			11'h467: data_out = 8'b01101000; // 7  ** *
			11'h468: data_out = 8'b01100000; // 8  **
			11'h469: data_out = 8'b01100000; // 9  **
			11'h46a: data_out = 8'b01100000; // a  **
			11'h46b: data_out = 8'b11110000; // b ****
			11'h46c: data_out = 8'b00000000; // c
			11'h46d: data_out = 8'b00000000; // d
			11'h46e: data_out = 8'b00000000; // e
			11'h46f: data_out = 8'b00000000; // f
			// code x47
			11'h470: data_out = 8'b00000000; // 0
			11'h471: data_out = 8'b00000000; // 1
			11'h472: data_out = 8'b00111100; // 2   ****
			11'h473: data_out = 8'b01100110; // 3  **  **
			11'h474: data_out = 8'b11000010; // 4 **    *
			11'h475: data_out = 8'b11000000; // 5 **
			11'h476: data_out = 8'b11000000; // 6 **
			11'h477: data_out = 8'b11011110; // 7 ** ****
			11'h478: data_out = 8'b11000110; // 8 **   **
			11'h479: data_out = 8'b11000110; // 9 **   **
			11'h47a: data_out = 8'b01100110; // a  **  **
			11'h47b: data_out = 8'b00111010; // b   *** *
			11'h47c: data_out = 8'b00000000; // c
			11'h47d: data_out = 8'b00000000; // d
			11'h47e: data_out = 8'b00000000; // e
			11'h47f: data_out = 8'b00000000; // f
			// code x48
			11'h480: data_out = 8'b00000000; // 0
			11'h481: data_out = 8'b00000000; // 1
			11'h482: data_out = 8'b11000110; // 2 **   **
			11'h483: data_out = 8'b11000110; // 3 **   **
			11'h484: data_out = 8'b11000110; // 4 **   **
			11'h485: data_out = 8'b11000110; // 5 **   **
			11'h486: data_out = 8'b11111110; // 6 *******
			11'h487: data_out = 8'b11000110; // 7 **   **
			11'h488: data_out = 8'b11000110; // 8 **   **
			11'h489: data_out = 8'b11000110; // 9 **   **
			11'h48a: data_out = 8'b11000110; // a **   **
			11'h48b: data_out = 8'b11000110; // b **   **
			11'h48c: data_out = 8'b00000000; // c
			11'h48d: data_out = 8'b00000000; // d
			11'h48e: data_out = 8'b00000000; // e
			11'h48f: data_out = 8'b00000000; // f
			// code x49
			11'h490: data_out = 8'b00000000; // 0
			11'h491: data_out = 8'b00000000; // 1
			11'h492: data_out = 8'b00111100; // 2   ****
			11'h493: data_out = 8'b00011000; // 3    **
			11'h494: data_out = 8'b00011000; // 4    **
			11'h495: data_out = 8'b00011000; // 5    **
			11'h496: data_out = 8'b00011000; // 6    **
			11'h497: data_out = 8'b00011000; // 7    **
			11'h498: data_out = 8'b00011000; // 8    **
			11'h499: data_out = 8'b00011000; // 9    **
			11'h49a: data_out = 8'b00011000; // a    **
			11'h49b: data_out = 8'b00111100; // b   ****
			11'h49c: data_out = 8'b00000000; // c
			11'h49d: data_out = 8'b00000000; // d
			11'h49e: data_out = 8'b00000000; // e
			11'h49f: data_out = 8'b00000000; // f
			// code x4a
			11'h4a0: data_out = 8'b00000000; // 0
			11'h4a1: data_out = 8'b00000000; // 1
			11'h4a2: data_out = 8'b00011110; // 2    ****
			11'h4a3: data_out = 8'b00001100; // 3     **
			11'h4a4: data_out = 8'b00001100; // 4     **
			11'h4a5: data_out = 8'b00001100; // 5     **
			11'h4a6: data_out = 8'b00001100; // 6     **
			11'h4a7: data_out = 8'b00001100; // 7     **
			11'h4a8: data_out = 8'b11001100; // 8 **  **
			11'h4a9: data_out = 8'b11001100; // 9 **  **
			11'h4aa: data_out = 8'b11001100; // a **  **
			11'h4ab: data_out = 8'b01111000; // b  ****
			11'h4ac: data_out = 8'b00000000; // c
			11'h4ad: data_out = 8'b00000000; // d
			11'h4ae: data_out = 8'b00000000; // e
			11'h4af: data_out = 8'b00000000; // f
			// code x4b
			11'h4b0: data_out = 8'b00000000; // 0
			11'h4b1: data_out = 8'b00000000; // 1
			11'h4b2: data_out = 8'b11100110; // 2 ***  **
			11'h4b3: data_out = 8'b01100110; // 3  **  **
			11'h4b4: data_out = 8'b01100110; // 4  **  **
			11'h4b5: data_out = 8'b01101100; // 5  ** **
			11'h4b6: data_out = 8'b01111000; // 6  ****
			11'h4b7: data_out = 8'b01111000; // 7  ****
			11'h4b8: data_out = 8'b01101100; // 8  ** **
			11'h4b9: data_out = 8'b01100110; // 9  **  **
			11'h4ba: data_out = 8'b01100110; // a  **  **
			11'h4bb: data_out = 8'b11100110; // b ***  **
			11'h4bc: data_out = 8'b00000000; // c
			11'h4bd: data_out = 8'b00000000; // d
			11'h4be: data_out = 8'b00000000; // e
			11'h4bf: data_out = 8'b00000000; // f
			// code x4c
			11'h4c0: data_out = 8'b00000000; // 0
			11'h4c1: data_out = 8'b00000000; // 1
			11'h4c2: data_out = 8'b11110000; // 2 ****
			11'h4c3: data_out = 8'b01100000; // 3  **
			11'h4c4: data_out = 8'b01100000; // 4  **
			11'h4c5: data_out = 8'b01100000; // 5  **
			11'h4c6: data_out = 8'b01100000; // 6  **
			11'h4c7: data_out = 8'b01100000; // 7  **
			11'h4c8: data_out = 8'b01100000; // 8  **
			11'h4c9: data_out = 8'b01100010; // 9  **   *
			11'h4ca: data_out = 8'b01100110; // a  **  **
			11'h4cb: data_out = 8'b11111110; // b *******
			11'h4cc: data_out = 8'b00000000; // c
			11'h4cd: data_out = 8'b00000000; // d
			11'h4ce: data_out = 8'b00000000; // e
			11'h4cf: data_out = 8'b00000000; // f
			// code x4d
			11'h4d0: data_out = 8'b00000000; // 0
			11'h4d1: data_out = 8'b00000000; // 1
			11'h4d2: data_out = 8'b11000011; // 2 **    **
			11'h4d3: data_out = 8'b11100111; // 3 ***  ***
			11'h4d4: data_out = 8'b11111111; // 4 ********
			11'h4d5: data_out = 8'b11111111; // 5 ********
			11'h4d6: data_out = 8'b11011011; // 6 ** ** **
			11'h4d7: data_out = 8'b11000011; // 7 **    **
			11'h4d8: data_out = 8'b11000011; // 8 **    **
			11'h4d9: data_out = 8'b11000011; // 9 **    **
			11'h4da: data_out = 8'b11000011; // a **    **
			11'h4db: data_out = 8'b11000011; // b **    **
			11'h4dc: data_out = 8'b00000000; // c
			11'h4dd: data_out = 8'b00000000; // d
			11'h4de: data_out = 8'b00000000; // e
			11'h4df: data_out = 8'b00000000; // f
			// code x4e
			11'h4e0: data_out = 8'b00000000; // 0
			11'h4e1: data_out = 8'b00000000; // 1
			11'h4e2: data_out = 8'b11000110; // 2 **   **
			11'h4e3: data_out = 8'b11100110; // 3 ***  **
			11'h4e4: data_out = 8'b11110110; // 4 **** **
			11'h4e5: data_out = 8'b11111110; // 5 *******
			11'h4e6: data_out = 8'b11011110; // 6 ** ****
			11'h4e7: data_out = 8'b11001110; // 7 **  ***
			11'h4e8: data_out = 8'b11000110; // 8 **   **
			11'h4e9: data_out = 8'b11000110; // 9 **   **
			11'h4ea: data_out = 8'b11000110; // a **   **
			11'h4eb: data_out = 8'b11000110; // b **   **
			11'h4ec: data_out = 8'b00000000; // c
			11'h4ed: data_out = 8'b00000000; // d
			11'h4ee: data_out = 8'b00000000; // e
			11'h4ef: data_out = 8'b00000000; // f
			// code x4f
			11'h4f0: data_out = 8'b00000000; // 0
			11'h4f1: data_out = 8'b00000000; // 1
			11'h4f2: data_out = 8'b01111100; // 2  *****
			11'h4f3: data_out = 8'b11000110; // 3 **   **
			11'h4f4: data_out = 8'b11000110; // 4 **   **
			11'h4f5: data_out = 8'b11000110; // 5 **   **
			11'h4f6: data_out = 8'b11000110; // 6 **   **
			11'h4f7: data_out = 8'b11000110; // 7 **   **
			11'h4f8: data_out = 8'b11000110; // 8 **   **
			11'h4f9: data_out = 8'b11000110; // 9 **   **
			11'h4fa: data_out = 8'b11000110; // a **   **
			11'h4fb: data_out = 8'b01111100; // b  *****
			11'h4fc: data_out = 8'b00000000; // c
			11'h4fd: data_out = 8'b00000000; // d
			11'h4fe: data_out = 8'b00000000; // e
			11'h4ff: data_out = 8'b00000000; // f
			// code x50
			11'h500: data_out = 8'b00000000; // 0
			11'h501: data_out = 8'b00000000; // 1
			11'h502: data_out = 8'b11111100; // 2 ******
			11'h503: data_out = 8'b01100110; // 3  **  **
			11'h504: data_out = 8'b01100110; // 4  **  **
			11'h505: data_out = 8'b01100110; // 5  **  **
			11'h506: data_out = 8'b01111100; // 6  *****
			11'h507: data_out = 8'b01100000; // 7  **
			11'h508: data_out = 8'b01100000; // 8  **
			11'h509: data_out = 8'b01100000; // 9  **
			11'h50a: data_out = 8'b01100000; // a  **
			11'h50b: data_out = 8'b11110000; // b ****
			11'h50c: data_out = 8'b00000000; // c
			11'h50d: data_out = 8'b00000000; // d
			11'h50e: data_out = 8'b00000000; // e
			11'h50f: data_out = 8'b00000000; // f
			// code x510
			11'h510: data_out = 8'b00000000; // 0
			11'h511: data_out = 8'b00000000; // 1
			11'h512: data_out = 8'b01111100; // 2  *****
			11'h513: data_out = 8'b11000110; // 3 **   **
			11'h514: data_out = 8'b11000110; // 4 **   **
			11'h515: data_out = 8'b11000110; // 5 **   **
			11'h516: data_out = 8'b11000110; // 6 **   **
			11'h517: data_out = 8'b11000110; // 7 **   **
			11'h518: data_out = 8'b11000110; // 8 **   **
			11'h519: data_out = 8'b11010110; // 9 ** * **
			11'h51a: data_out = 8'b11011110; // a ** ****
			11'h51b: data_out = 8'b01111100; // b  *****
			11'h51c: data_out = 8'b00001100; // c     **
			11'h51d: data_out = 8'b00001110; // d     ***
			11'h51e: data_out = 8'b00000000; // e
			11'h51f: data_out = 8'b00000000; // f
			// code x52
			11'h520: data_out = 8'b00000000; // 0
			11'h521: data_out = 8'b00000000; // 1
			11'h522: data_out = 8'b11111100; // 2 ******
			11'h523: data_out = 8'b01100110; // 3  **  **
			11'h524: data_out = 8'b01100110; // 4  **  **
			11'h525: data_out = 8'b01100110; // 5  **  **
			11'h526: data_out = 8'b01111100; // 6  *****
			11'h527: data_out = 8'b01101100; // 7  ** **
			11'h528: data_out = 8'b01100110; // 8  **  **
			11'h529: data_out = 8'b01100110; // 9  **  **
			11'h52a: data_out = 8'b01100110; // a  **  **
			11'h52b: data_out = 8'b11100110; // b ***  **
			11'h52c: data_out = 8'b00000000; // c
			11'h52d: data_out = 8'b00000000; // d
			11'h52e: data_out = 8'b00000000; // e
			11'h52f: data_out = 8'b00000000; // f
			// code x53
			11'h530: data_out = 8'b00000000; // 0
			11'h531: data_out = 8'b00000000; // 1
			11'h532: data_out = 8'b01111100; // 2  *****
			11'h533: data_out = 8'b11000110; // 3 **   **
			11'h534: data_out = 8'b11000110; // 4 **   **
			11'h535: data_out = 8'b01100000; // 5  **
			11'h536: data_out = 8'b00111000; // 6   ***
			11'h537: data_out = 8'b00001100; // 7     **
			11'h538: data_out = 8'b00000110; // 8      **
			11'h539: data_out = 8'b11000110; // 9 **   **
			11'h53a: data_out = 8'b11000110; // a **   **
			11'h53b: data_out = 8'b01111100; // b  *****
			11'h53c: data_out = 8'b00000000; // c
			11'h53d: data_out = 8'b00000000; // d
			11'h53e: data_out = 8'b00000000; // e
			11'h53f: data_out = 8'b00000000; // f
			// code x54
			11'h540: data_out = 8'b00000000; // 0
			11'h541: data_out = 8'b00000000; // 1
			11'h542: data_out = 8'b11111111; // 2 ********
			11'h543: data_out = 8'b11011011; // 3 ** ** **
			11'h544: data_out = 8'b10011001; // 4 *  **  *
			11'h545: data_out = 8'b00011000; // 5    **
			11'h546: data_out = 8'b00011000; // 6    **
			11'h547: data_out = 8'b00011000; // 7    **
			11'h548: data_out = 8'b00011000; // 8    **
			11'h549: data_out = 8'b00011000; // 9    **
			11'h54a: data_out = 8'b00011000; // a    **
			11'h54b: data_out = 8'b00111100; // b   ****
			11'h54c: data_out = 8'b00000000; // c
			11'h54d: data_out = 8'b00000000; // d
			11'h54e: data_out = 8'b00000000; // e
			11'h54f: data_out = 8'b00000000; // f
			// code x55
			11'h550: data_out = 8'b00000000; // 0
			11'h551: data_out = 8'b00000000; // 1
			11'h552: data_out = 8'b11000110; // 2 **   **
			11'h553: data_out = 8'b11000110; // 3 **   **
			11'h554: data_out = 8'b11000110; // 4 **   **
			11'h555: data_out = 8'b11000110; // 5 **   **
			11'h556: data_out = 8'b11000110; // 6 **   **
			11'h557: data_out = 8'b11000110; // 7 **   **
			11'h558: data_out = 8'b11000110; // 8 **   **
			11'h559: data_out = 8'b11000110; // 9 **   **
			11'h55a: data_out = 8'b11000110; // a **   **
			11'h55b: data_out = 8'b01111100; // b  *****
			11'h55c: data_out = 8'b00000000; // c
			11'h55d: data_out = 8'b00000000; // d
			11'h55e: data_out = 8'b00000000; // e
			11'h55f: data_out = 8'b00000000; // f
			// code x56
			11'h560: data_out = 8'b00000000; // 0
			11'h561: data_out = 8'b00000000; // 1
			11'h562: data_out = 8'b11000011; // 2 **    **
			11'h563: data_out = 8'b11000011; // 3 **    **
			11'h564: data_out = 8'b11000011; // 4 **    **
			11'h565: data_out = 8'b11000011; // 5 **    **
			11'h566: data_out = 8'b11000011; // 6 **    **
			11'h567: data_out = 8'b11000011; // 7 **    **
			11'h568: data_out = 8'b11000011; // 8 **    **
			11'h569: data_out = 8'b01100110; // 9  **  **
			11'h56a: data_out = 8'b00111100; // a   ****
			11'h56b: data_out = 8'b00011000; // b    **
			11'h56c: data_out = 8'b00000000; // c
			11'h56d: data_out = 8'b00000000; // d
			11'h56e: data_out = 8'b00000000; // e
			11'h56f: data_out = 8'b00000000; // f
			// code x57
			11'h570: data_out = 8'b00000000; // 0
			11'h571: data_out = 8'b00000000; // 1
			11'h572: data_out = 8'b11000011; // 2 **    **
			11'h573: data_out = 8'b11000011; // 3 **    **
			11'h574: data_out = 8'b11000011; // 4 **    **
			11'h575: data_out = 8'b11000011; // 5 **    **
			11'h576: data_out = 8'b11000011; // 6 **    **
			11'h577: data_out = 8'b11011011; // 7 ** ** **
			11'h578: data_out = 8'b11011011; // 8 ** ** **
			11'h579: data_out = 8'b11111111; // 9 ********
			11'h57a: data_out = 8'b01100110; // a  **  **
			11'h57b: data_out = 8'b01100110; // b  **  **
			11'h57c: data_out = 8'b00000000; // c
			11'h57d: data_out = 8'b00000000; // d
			11'h57e: data_out = 8'b00000000; // e
			11'h57f: data_out = 8'b00000000; // f

			// code x58
			11'h580: data_out = 8'b00000000; // 0
			11'h581: data_out = 8'b00000000; // 1
			11'h582: data_out = 8'b11000011; // 2 **    **
			11'h583: data_out = 8'b11000011; // 3 **    **
			11'h584: data_out = 8'b01100110; // 4  **  **
			11'h585: data_out = 8'b00111100; // 5   ****
			11'h586: data_out = 8'b00011000; // 6    **
			11'h587: data_out = 8'b00011000; // 7    **
			11'h588: data_out = 8'b00111100; // 8   ****
			11'h589: data_out = 8'b01100110; // 9  **  **
			11'h58a: data_out = 8'b11000011; // a **    **
			11'h58b: data_out = 8'b11000011; // b **    **
			11'h58c: data_out = 8'b00000000; // c
			11'h58d: data_out = 8'b00000000; // d
			11'h58e: data_out = 8'b00000000; // e
			11'h58f: data_out = 8'b00000000; // f
			// code x59
			11'h590: data_out = 8'b00000000; // 0
			11'h591: data_out = 8'b00000000; // 1
			11'h592: data_out = 8'b11000011; // 2 **    **
			11'h593: data_out = 8'b11000011; // 3 **    **
			11'h594: data_out = 8'b11000011; // 4 **    **
			11'h595: data_out = 8'b01100110; // 5  **  **
			11'h596: data_out = 8'b00111100; // 6   ****
			11'h597: data_out = 8'b00011000; // 7    **
			11'h598: data_out = 8'b00011000; // 8    **
			11'h599: data_out = 8'b00011000; // 9    **
			11'h59a: data_out = 8'b00011000; // a    **
			11'h59b: data_out = 8'b00111100; // b   ****
			11'h59c: data_out = 8'b00000000; // c
			11'h59d: data_out = 8'b00000000; // d
			11'h59e: data_out = 8'b00000000; // e
			11'h59f: data_out = 8'b00000000; // f
			// code x5a
			11'h5a0: data_out = 8'b00000000; // 0
			11'h5a1: data_out = 8'b00000000; // 1
			11'h5a2: data_out = 8'b11111111; // 2 ********
			11'h5a3: data_out = 8'b11000011; // 3 **    **
			11'h5a4: data_out = 8'b10000110; // 4 *    **
			11'h5a5: data_out = 8'b00001100; // 5     **
			11'h5a6: data_out = 8'b00011000; // 6    **
			11'h5a7: data_out = 8'b00110000; // 7   **
			11'h5a8: data_out = 8'b01100000; // 8  **
			11'h5a9: data_out = 8'b11000001; // 9 **     *
			11'h5aa: data_out = 8'b11000011; // a **    **
			11'h5ab: data_out = 8'b11111111; // b ********
			11'h5ac: data_out = 8'b00000000; // c
			11'h5ad: data_out = 8'b00000000; // d
			11'h5ae: data_out = 8'b00000000; // e
			11'h5af: data_out = 8'b00000000; // f
			// code x5b
			11'h5b0: data_out = 8'b00000000; // 0
			11'h5b1: data_out = 8'b00000000; // 1
			11'h5b2: data_out = 8'b00111100; // 2   ****
			11'h5b3: data_out = 8'b00110000; // 3   **
			11'h5b4: data_out = 8'b00110000; // 4   **
			11'h5b5: data_out = 8'b00110000; // 5   **
			11'h5b6: data_out = 8'b00110000; // 6   **
			11'h5b7: data_out = 8'b00110000; // 7   **
			11'h5b8: data_out = 8'b00110000; // 8   **
			11'h5b9: data_out = 8'b00110000; // 9   **
			11'h5ba: data_out = 8'b00110000; // a   **
			11'h5bb: data_out = 8'b00111100; // b   ****
			11'h5bc: data_out = 8'b00000000; // c
			11'h5bd: data_out = 8'b00000000; // d
			11'h5be: data_out = 8'b00000000; // e
			11'h5bf: data_out = 8'b00000000; // f
			// code x5c
			11'h5c0: data_out = 8'b00000000; // 0
			11'h5c1: data_out = 8'b00000000; // 1
			11'h5c2: data_out = 8'b00000000; // 2
			11'h5c3: data_out = 8'b10000000; // 3 *
			11'h5c4: data_out = 8'b11000000; // 4 **
			11'h5c5: data_out = 8'b11100000; // 5 ***
			11'h5c6: data_out = 8'b01110000; // 6  ***
			11'h5c7: data_out = 8'b00111000; // 7   ***
			11'h5c8: data_out = 8'b00011100; // 8    ***
			11'h5c9: data_out = 8'b00001110; // 9     ***
			11'h5ca: data_out = 8'b00000110; // a      **
			11'h5cb: data_out = 8'b00000010; // b       *
			11'h5cc: data_out = 8'b00000000; // c
			11'h5cd: data_out = 8'b00000000; // d
			11'h5ce: data_out = 8'b00000000; // e
			11'h5cf: data_out = 8'b00000000; // f
			// code x5d
			11'h5d0: data_out = 8'b00000000; // 0
			11'h5d1: data_out = 8'b00000000; // 1
			11'h5d2: data_out = 8'b00111100; // 2   ****
			11'h5d3: data_out = 8'b00001100; // 3     **
			11'h5d4: data_out = 8'b00001100; // 4     **
			11'h5d5: data_out = 8'b00001100; // 5     **
			11'h5d6: data_out = 8'b00001100; // 6     **
			11'h5d7: data_out = 8'b00001100; // 7     **
			11'h5d8: data_out = 8'b00001100; // 8     **
			11'h5d9: data_out = 8'b00001100; // 9     **
			11'h5da: data_out = 8'b00001100; // a     **
			11'h5db: data_out = 8'b00111100; // b   ****
			11'h5dc: data_out = 8'b00000000; // c
			11'h5dd: data_out = 8'b00000000; // d
			11'h5de: data_out = 8'b00000000; // e
			11'h5df: data_out = 8'b00000000; // f
			// code x5e
			11'h5e0: data_out = 8'b00010000; // 0    *
			11'h5e1: data_out = 8'b00111000; // 1   ***
			11'h5e2: data_out = 8'b01101100; // 2  ** **
			11'h5e3: data_out = 8'b11000110; // 3 **   **
			11'h5e4: data_out = 8'b00000000; // 4
			11'h5e5: data_out = 8'b00000000; // 5
			11'h5e6: data_out = 8'b00000000; // 6
			11'h5e7: data_out = 8'b00000000; // 7
			11'h5e8: data_out = 8'b00000000; // 8
			11'h5e9: data_out = 8'b00000000; // 9
			11'h5ea: data_out = 8'b00000000; // a
			11'h5eb: data_out = 8'b00000000; // b
			11'h5ec: data_out = 8'b00000000; // c
			11'h5ed: data_out = 8'b00000000; // d
			11'h5ee: data_out = 8'b00000000; // e
			11'h5ef: data_out = 8'b00000000; // f
			// code x5f
			11'h5f0: data_out = 8'b00000000; // 0
			11'h5f1: data_out = 8'b00000000; // 1
			11'h5f2: data_out = 8'b00000000; // 2
			11'h5f3: data_out = 8'b00000000; // 3
			11'h5f4: data_out = 8'b00000000; // 4
			11'h5f5: data_out = 8'b00000000; // 5
			11'h5f6: data_out = 8'b00000000; // 6
			11'h5f7: data_out = 8'b00000000; // 7
			11'h5f8: data_out = 8'b00000000; // 8
			11'h5f9: data_out = 8'b00000000; // 9
			11'h5fa: data_out = 8'b00000000; // a
			11'h5fb: data_out = 8'b00000000; // b
			11'h5fc: data_out = 8'b00000000; // c
			11'h5fd: data_out = 8'b11111111; // d ********
			11'h5fe: data_out = 8'b00000000; // e
			11'h5ff: data_out = 8'b00000000; // f
			// code x60
			11'h600: data_out = 8'b00110000; // 0   **
			11'h601: data_out = 8'b00110000; // 1   **
			11'h602: data_out = 8'b00011000; // 2    **
			11'h603: data_out = 8'b00000000; // 3
			11'h604: data_out = 8'b00000000; // 4
			11'h605: data_out = 8'b00000000; // 5
			11'h606: data_out = 8'b00000000; // 6
			11'h607: data_out = 8'b00000000; // 7
			11'h608: data_out = 8'b00000000; // 8
			11'h609: data_out = 8'b00000000; // 9
			11'h60a: data_out = 8'b00000000; // a
			11'h60b: data_out = 8'b00000000; // b
			11'h60c: data_out = 8'b00000000; // c
			11'h60d: data_out = 8'b00000000; // d
			11'h60e: data_out = 8'b00000000; // e
			11'h60f: data_out = 8'b00000000; // f
			// code x61
			11'h610: data_out = 8'b00000000; // 0
			11'h611: data_out = 8'b00000000; // 1
			11'h612: data_out = 8'b00000000; // 2
			11'h613: data_out = 8'b00000000; // 3
			11'h614: data_out = 8'b00000000; // 4
			11'h615: data_out = 8'b01111000; // 5  ****
			11'h616: data_out = 8'b00001100; // 6     **
			11'h617: data_out = 8'b01111100; // 7  *****
			11'h618: data_out = 8'b11001100; // 8 **  **
			11'h619: data_out = 8'b11001100; // 9 **  **
			11'h61a: data_out = 8'b11001100; // a **  **
			11'h61b: data_out = 8'b01110110; // b  *** **
			11'h61c: data_out = 8'b00000000; // c
			11'h61d: data_out = 8'b00000000; // d
			11'h61e: data_out = 8'b00000000; // e
			11'h61f: data_out = 8'b00000000; // f
			// code x62
			11'h620: data_out = 8'b00000000; // 0
			11'h621: data_out = 8'b00000000; // 1
			11'h622: data_out = 8'b11100000; // 2  ***
			11'h623: data_out = 8'b01100000; // 3   **
			11'h624: data_out = 8'b01100000; // 4   **
			11'h625: data_out = 8'b01111000; // 5   ****
			11'h626: data_out = 8'b01101100; // 6   ** **
			11'h627: data_out = 8'b01100110; // 7   **  **
			11'h628: data_out = 8'b01100110; // 8   **  **
			11'h629: data_out = 8'b01100110; // 9   **  **
			11'h62a: data_out = 8'b01100110; // a   **  **
			11'h62b: data_out = 8'b01111100; // b   *****
			11'h62c: data_out = 8'b00000000; // c
			11'h62d: data_out = 8'b00000000; // d
			11'h62e: data_out = 8'b00000000; // e
			11'h62f: data_out = 8'b00000000; // f
			// code x63
			11'h630: data_out = 8'b00000000; // 0
			11'h631: data_out = 8'b00000000; // 1
			11'h632: data_out = 8'b00000000; // 2
			11'h633: data_out = 8'b00000000; // 3
			11'h634: data_out = 8'b00000000; // 4
			11'h635: data_out = 8'b01111100; // 5  *****
			11'h636: data_out = 8'b11000110; // 6 **   **
			11'h637: data_out = 8'b11000000; // 7 **
			11'h638: data_out = 8'b11000000; // 8 **
			11'h639: data_out = 8'b11000000; // 9 **
			11'h63a: data_out = 8'b11000110; // a **   **
			11'h63b: data_out = 8'b01111100; // b  *****
			11'h63c: data_out = 8'b00000000; // c
			11'h63d: data_out = 8'b00000000; // d
			11'h63e: data_out = 8'b00000000; // e
			11'h63f: data_out = 8'b00000000; // f
			// code x64
			11'h640: data_out = 8'b00000000; // 0
			11'h641: data_out = 8'b00000000; // 1
			11'h642: data_out = 8'b00011100; // 2    ***
			11'h643: data_out = 8'b00001100; // 3     **
			11'h644: data_out = 8'b00001100; // 4     **
			11'h645: data_out = 8'b00111100; // 5   ****
			11'h646: data_out = 8'b01101100; // 6  ** **
			11'h647: data_out = 8'b11001100; // 7 **  **
			11'h648: data_out = 8'b11001100; // 8 **  **
			11'h649: data_out = 8'b11001100; // 9 **  **
			11'h64a: data_out = 8'b11001100; // a **  **
			11'h64b: data_out = 8'b01110110; // b  *** **
			11'h64c: data_out = 8'b00000000; // c
			11'h64d: data_out = 8'b00000000; // d
			11'h64e: data_out = 8'b00000000; // e
			11'h64f: data_out = 8'b00000000; // f
			// code x65
			11'h650: data_out = 8'b00000000; // 0
			11'h651: data_out = 8'b00000000; // 1
			11'h652: data_out = 8'b00000000; // 2
			11'h653: data_out = 8'b00000000; // 3
			11'h654: data_out = 8'b00000000; // 4
			11'h655: data_out = 8'b01111100; // 5  *****
			11'h656: data_out = 8'b11000110; // 6 **   **
			11'h657: data_out = 8'b11111110; // 7 *******
			11'h658: data_out = 8'b11000000; // 8 **
			11'h659: data_out = 8'b11000000; // 9 **
			11'h65a: data_out = 8'b11000110; // a **   **
			11'h65b: data_out = 8'b01111100; // b  *****
			11'h65c: data_out = 8'b00000000; // c
			11'h65d: data_out = 8'b00000000; // d
			11'h65e: data_out = 8'b00000000; // e
			11'h65f: data_out = 8'b00000000; // f
			// code x66
			11'h660: data_out = 8'b00000000; // 0
			11'h661: data_out = 8'b00000000; // 1
			11'h662: data_out = 8'b00111000; // 2   ***
			11'h663: data_out = 8'b01101100; // 3  ** **
			11'h664: data_out = 8'b01100100; // 4  **  *
			11'h665: data_out = 8'b01100000; // 5  **
			11'h666: data_out = 8'b11110000; // 6 ****
			11'h667: data_out = 8'b01100000; // 7  **
			11'h668: data_out = 8'b01100000; // 8  **
			11'h669: data_out = 8'b01100000; // 9  **
			11'h66a: data_out = 8'b01100000; // a  **
			11'h66b: data_out = 8'b11110000; // b ****
			11'h66c: data_out = 8'b00000000; // c
			11'h66d: data_out = 8'b00000000; // d
			11'h66e: data_out = 8'b00000000; // e
			11'h66f: data_out = 8'b00000000; // f
			// code x67
			11'h670: data_out = 8'b00000000; // 0
			11'h671: data_out = 8'b00000000; // 1
			11'h672: data_out = 8'b00000000; // 2
			11'h673: data_out = 8'b00000000; // 3
			11'h674: data_out = 8'b00000000; // 4
			11'h675: data_out = 8'b01110110; // 5  *** **
			11'h676: data_out = 8'b11001100; // 6 **  **
			11'h677: data_out = 8'b11001100; // 7 **  **
			11'h678: data_out = 8'b11001100; // 8 **  **
			11'h679: data_out = 8'b11001100; // 9 **  **
			11'h67a: data_out = 8'b11001100; // a **  **
			11'h67b: data_out = 8'b01111100; // b  *****
			11'h67c: data_out = 8'b00001100; // c     **
			11'h67d: data_out = 8'b11001100; // d **  **
			11'h67e: data_out = 8'b01111000; // e  ****
			11'h67f: data_out = 8'b00000000; // f
			// code x68
			11'h680: data_out = 8'b00000000; // 0
			11'h681: data_out = 8'b00000000; // 1
			11'h682: data_out = 8'b11100000; // 2 ***
			11'h683: data_out = 8'b01100000; // 3  **
			11'h684: data_out = 8'b01100000; // 4  **
			11'h685: data_out = 8'b01101100; // 5  ** **
			11'h686: data_out = 8'b01110110; // 6  *** **
			11'h687: data_out = 8'b01100110; // 7  **  **
			11'h688: data_out = 8'b01100110; // 8  **  **
			11'h689: data_out = 8'b01100110; // 9  **  **
			11'h68a: data_out = 8'b01100110; // a  **  **
			11'h68b: data_out = 8'b11100110; // b ***  **
			11'h68c: data_out = 8'b00000000; // c
			11'h68d: data_out = 8'b00000000; // d
			11'h68e: data_out = 8'b00000000; // e
			11'h68f: data_out = 8'b00000000; // f
			// code x69
			11'h690: data_out = 8'b00000000; // 0
			11'h691: data_out = 8'b00000000; // 1
			11'h692: data_out = 8'b00011000; // 2    **
			11'h693: data_out = 8'b00011000; // 3    **
			11'h694: data_out = 8'b00000000; // 4
			11'h695: data_out = 8'b00111000; // 5   ***
			11'h696: data_out = 8'b00011000; // 6    **
			11'h697: data_out = 8'b00011000; // 7    **
			11'h698: data_out = 8'b00011000; // 8    **
			11'h699: data_out = 8'b00011000; // 9    **
			11'h69a: data_out = 8'b00011000; // a    **
			11'h69b: data_out = 8'b00111100; // b   ****
			11'h69c: data_out = 8'b00000000; // c
			11'h69d: data_out = 8'b00000000; // d
			11'h69e: data_out = 8'b00000000; // e
			11'h69f: data_out = 8'b00000000; // f
			// code x6a
			11'h6a0: data_out = 8'b00000000; // 0
			11'h6a1: data_out = 8'b00000000; // 1
			11'h6a2: data_out = 8'b00000110; // 2      **
			11'h6a3: data_out = 8'b00000110; // 3      **
			11'h6a4: data_out = 8'b00000000; // 4
			11'h6a5: data_out = 8'b00001110; // 5     ***
			11'h6a6: data_out = 8'b00000110; // 6      **
			11'h6a7: data_out = 8'b00000110; // 7      **
			11'h6a8: data_out = 8'b00000110; // 8      **
			11'h6a9: data_out = 8'b00000110; // 9      **
			11'h6aa: data_out = 8'b00000110; // a      **
			11'h6ab: data_out = 8'b00000110; // b      **
			11'h6ac: data_out = 8'b01100110; // c  **  **
			11'h6ad: data_out = 8'b01100110; // d  **  **
			11'h6ae: data_out = 8'b00111100; // e   ****
			11'h6af: data_out = 8'b00000000; // f
			// code x6b
			11'h6b0: data_out = 8'b00000000; // 0
			11'h6b1: data_out = 8'b00000000; // 1
			11'h6b2: data_out = 8'b11100000; // 2 ***
			11'h6b3: data_out = 8'b01100000; // 3  **
			11'h6b4: data_out = 8'b01100000; // 4  **
			11'h6b5: data_out = 8'b01100110; // 5  **  **
			11'h6b6: data_out = 8'b01101100; // 6  ** **
			11'h6b7: data_out = 8'b01111000; // 7  ****
			11'h6b8: data_out = 8'b01111000; // 8  ****
			11'h6b9: data_out = 8'b01101100; // 9  ** **
			11'h6ba: data_out = 8'b01100110; // a  **  **
			11'h6bb: data_out = 8'b11100110; // b ***  **
			11'h6bc: data_out = 8'b00000000; // c
			11'h6bd: data_out = 8'b00000000; // d
			11'h6be: data_out = 8'b00000000; // e
			11'h6bf: data_out = 8'b00000000; // f
			// code x6c
			11'h6c0: data_out = 8'b00000000; // 0
			11'h6c1: data_out = 8'b00000000; // 1
			11'h6c2: data_out = 8'b00111000; // 2   ***
			11'h6c3: data_out = 8'b00011000; // 3    **
			11'h6c4: data_out = 8'b00011000; // 4    **
			11'h6c5: data_out = 8'b00011000; // 5    **
			11'h6c6: data_out = 8'b00011000; // 6    **
			11'h6c7: data_out = 8'b00011000; // 7    **
			11'h6c8: data_out = 8'b00011000; // 8    **
			11'h6c9: data_out = 8'b00011000; // 9    **
			11'h6ca: data_out = 8'b00011000; // a    **
			11'h6cb: data_out = 8'b00111100; // b   ****
			11'h6cc: data_out = 8'b00000000; // c
			11'h6cd: data_out = 8'b00000000; // d
			11'h6ce: data_out = 8'b00000000; // e
			11'h6cf: data_out = 8'b00000000; // f
			// code x6d
			11'h6d0: data_out = 8'b00000000; // 0
			11'h6d1: data_out = 8'b00000000; // 1
			11'h6d2: data_out = 8'b00000000; // 2
			11'h6d3: data_out = 8'b00000000; // 3
			11'h6d4: data_out = 8'b00000000; // 4
			11'h6d5: data_out = 8'b11100110; // 5 ***  **
			11'h6d6: data_out = 8'b11111111; // 6 ********
			11'h6d7: data_out = 8'b11011011; // 7 ** ** **
			11'h6d8: data_out = 8'b11011011; // 8 ** ** **
			11'h6d9: data_out = 8'b11011011; // 9 ** ** **
			11'h6da: data_out = 8'b11011011; // a ** ** **
			11'h6db: data_out = 8'b11011011; // b ** ** **
			11'h6dc: data_out = 8'b00000000; // c
			11'h6dd: data_out = 8'b00000000; // d
			11'h6de: data_out = 8'b00000000; // e
			11'h6df: data_out = 8'b00000000; // f
			// code x6e
			11'h6e0: data_out = 8'b00000000; // 0
			11'h6e1: data_out = 8'b00000000; // 1
			11'h6e2: data_out = 8'b00000000; // 2
			11'h6e3: data_out = 8'b00000000; // 3
			11'h6e4: data_out = 8'b00000000; // 4
			11'h6e5: data_out = 8'b11011100; // 5 ** ***
			11'h6e6: data_out = 8'b01100110; // 6  **  **
			11'h6e7: data_out = 8'b01100110; // 7  **  **
			11'h6e8: data_out = 8'b01100110; // 8  **  **
			11'h6e9: data_out = 8'b01100110; // 9  **  **
			11'h6ea: data_out = 8'b01100110; // a  **  **
			11'h6eb: data_out = 8'b01100110; // b  **  **
			11'h6ec: data_out = 8'b00000000; // c
			11'h6ed: data_out = 8'b00000000; // d
			11'h6ee: data_out = 8'b00000000; // e
			11'h6ef: data_out = 8'b00000000; // f
			// code x6f
			11'h6f0: data_out = 8'b00000000; // 0
			11'h6f1: data_out = 8'b00000000; // 1
			11'h6f2: data_out = 8'b00000000; // 2
			11'h6f3: data_out = 8'b00000000; // 3
			11'h6f4: data_out = 8'b00000000; // 4
			11'h6f5: data_out = 8'b01111100; // 5  *****
			11'h6f6: data_out = 8'b11000110; // 6 **   **
			11'h6f7: data_out = 8'b11000110; // 7 **   **
			11'h6f8: data_out = 8'b11000110; // 8 **   **
			11'h6f9: data_out = 8'b11000110; // 9 **   **
			11'h6fa: data_out = 8'b11000110; // a **   **
			11'h6fb: data_out = 8'b01111100; // b  *****
			11'h6fc: data_out = 8'b00000000; // c
			11'h6fd: data_out = 8'b00000000; // d
			11'h6fe: data_out = 8'b00000000; // e
			11'h6ff: data_out = 8'b00000000; // f
			// code x70
			11'h700: data_out = 8'b00000000; // 0
			11'h701: data_out = 8'b00000000; // 1
			11'h702: data_out = 8'b00000000; // 2
			11'h703: data_out = 8'b00000000; // 3
			11'h704: data_out = 8'b00000000; // 4
			11'h705: data_out = 8'b11011100; // 5 ** ***
			11'h706: data_out = 8'b01100110; // 6  **  **
			11'h707: data_out = 8'b01100110; // 7  **  **
			11'h708: data_out = 8'b01100110; // 8  **  **
			11'h709: data_out = 8'b01100110; // 9  **  **
			11'h70a: data_out = 8'b01100110; // a  **  **
			11'h70b: data_out = 8'b01111100; // b  *****
			11'h70c: data_out = 8'b01100000; // c  **
			11'h70d: data_out = 8'b01100000; // d  **
			11'h70e: data_out = 8'b11110000; // e ****
			11'h70f: data_out = 8'b00000000; // f
			// code x71
			11'h710: data_out = 8'b00000000; // 0
			11'h711: data_out = 8'b00000000; // 1
			11'h712: data_out = 8'b00000000; // 2
			11'h713: data_out = 8'b00000000; // 3
			11'h714: data_out = 8'b00000000; // 4
			11'h715: data_out = 8'b01110110; // 5  *** **
			11'h716: data_out = 8'b11001100; // 6 **  **
			11'h717: data_out = 8'b11001100; // 7 **  **
			11'h718: data_out = 8'b11001100; // 8 **  **
			11'h719: data_out = 8'b11001100; // 9 **  **
			11'h71a: data_out = 8'b11001100; // a **  **
			11'h71b: data_out = 8'b01111100; // b  *****
			11'h71c: data_out = 8'b00001100; // c     **
			11'h71d: data_out = 8'b00001100; // d     **
			11'h71e: data_out = 8'b00011110; // e    ****
			11'h71f: data_out = 8'b00000000; // f
			// code x72
			11'h720: data_out = 8'b00000000; // 0
			11'h721: data_out = 8'b00000000; // 1
			11'h722: data_out = 8'b00000000; // 2
			11'h723: data_out = 8'b00000000; // 3
			11'h724: data_out = 8'b00000000; // 4
			11'h725: data_out = 8'b11011100; // 5 ** ***
			11'h726: data_out = 8'b01110110; // 6  *** **
			11'h727: data_out = 8'b01100110; // 7  **  **
			11'h728: data_out = 8'b01100000; // 8  **
			11'h729: data_out = 8'b01100000; // 9  **
			11'h72a: data_out = 8'b01100000; // a  **
			11'h72b: data_out = 8'b11110000; // b ****
			11'h72c: data_out = 8'b00000000; // c
			11'h72d: data_out = 8'b00000000; // d
			11'h72e: data_out = 8'b00000000; // e
			11'h72f: data_out = 8'b00000000; // f
			// code x73
			11'h730: data_out = 8'b00000000; // 0
			11'h731: data_out = 8'b00000000; // 1
			11'h732: data_out = 8'b00000000; // 2
			11'h733: data_out = 8'b00000000; // 3
			11'h734: data_out = 8'b00000000; // 4
			11'h735: data_out = 8'b01111100; // 5  *****
			11'h736: data_out = 8'b11000110; // 6 **   **
			11'h737: data_out = 8'b01100000; // 7  **
			11'h738: data_out = 8'b00111000; // 8   ***
			11'h739: data_out = 8'b00001100; // 9     **
			11'h73a: data_out = 8'b11000110; // a **   **
			11'h73b: data_out = 8'b01111100; // b  *****
			11'h73c: data_out = 8'b00000000; // c
			11'h73d: data_out = 8'b00000000; // d
			11'h73e: data_out = 8'b00000000; // e
			11'h73f: data_out = 8'b00000000; // f
			// code x74
			11'h740: data_out = 8'b00000000; // 0
			11'h741: data_out = 8'b00000000; // 1
			11'h742: data_out = 8'b00010000; // 2    *
			11'h743: data_out = 8'b00110000; // 3   **
			11'h744: data_out = 8'b00110000; // 4   **
			11'h745: data_out = 8'b11111100; // 5 ******
			11'h746: data_out = 8'b00110000; // 6   **
			11'h747: data_out = 8'b00110000; // 7   **
			11'h748: data_out = 8'b00110000; // 8   **
			11'h749: data_out = 8'b00110000; // 9   **
			11'h74a: data_out = 8'b00110110; // a   ** **
			11'h74b: data_out = 8'b00011100; // b    ***
			11'h74c: data_out = 8'b00000000; // c
			11'h74d: data_out = 8'b00000000; // d
			11'h74e: data_out = 8'b00000000; // e
			11'h74f: data_out = 8'b00000000; // f
			// code x75
			11'h750: data_out = 8'b00000000; // 0
			11'h751: data_out = 8'b00000000; // 1
			11'h752: data_out = 8'b00000000; // 2
			11'h753: data_out = 8'b00000000; // 3
			11'h754: data_out = 8'b00000000; // 4
			11'h755: data_out = 8'b11001100; // 5 **  **
			11'h756: data_out = 8'b11001100; // 6 **  **
			11'h757: data_out = 8'b11001100; // 7 **  **
			11'h758: data_out = 8'b11001100; // 8 **  **
			11'h759: data_out = 8'b11001100; // 9 **  **
			11'h75a: data_out = 8'b11001100; // a **  **
			11'h75b: data_out = 8'b01110110; // b  *** **
			11'h75c: data_out = 8'b00000000; // c
			11'h75d: data_out = 8'b00000000; // d
			11'h75e: data_out = 8'b00000000; // e
			11'h75f: data_out = 8'b00000000; // f
			// code x76
			11'h760: data_out = 8'b00000000; // 0
			11'h761: data_out = 8'b00000000; // 1
			11'h762: data_out = 8'b00000000; // 2
			11'h763: data_out = 8'b00000000; // 3
			11'h764: data_out = 8'b00000000; // 4
			11'h765: data_out = 8'b11000011; // 5 **    **
			11'h766: data_out = 8'b11000011; // 6 **    **
			11'h767: data_out = 8'b11000011; // 7 **    **
			11'h768: data_out = 8'b11000011; // 8 **    **
			11'h769: data_out = 8'b01100110; // 9  **  **
			11'h76a: data_out = 8'b00111100; // a   ****
			11'h76b: data_out = 8'b00011000; // b    **
			11'h76c: data_out = 8'b00000000; // c
			11'h76d: data_out = 8'b00000000; // d
			11'h76e: data_out = 8'b00000000; // e
			11'h76f: data_out = 8'b00000000; // f
			// code x77
			11'h770: data_out = 8'b00000000; // 0
			11'h771: data_out = 8'b00000000; // 1
			11'h772: data_out = 8'b00000000; // 2
			11'h773: data_out = 8'b00000000; // 3
			11'h774: data_out = 8'b00000000; // 4
			11'h775: data_out = 8'b11000011; // 5 **    **
			11'h776: data_out = 8'b11000011; // 6 **    **
			11'h777: data_out = 8'b11000011; // 7 **    **
			11'h778: data_out = 8'b11011011; // 8 ** ** **
			11'h779: data_out = 8'b11011011; // 9 ** ** **
			11'h77a: data_out = 8'b11111111; // a ********
			11'h77b: data_out = 8'b01100110; // b  **  **
			11'h77c: data_out = 8'b00000000; // c
			11'h77d: data_out = 8'b00000000; // d
			11'h77e: data_out = 8'b00000000; // e
			11'h77f: data_out = 8'b00000000; // f
			// code x78
			11'h780: data_out = 8'b00000000; // 0
			11'h781: data_out = 8'b00000000; // 1
			11'h782: data_out = 8'b00000000; // 2
			11'h783: data_out = 8'b00000000; // 3
			11'h784: data_out = 8'b00000000; // 4
			11'h785: data_out = 8'b11000011; // 5 **    **
			11'h786: data_out = 8'b01100110; // 6  **  **
			11'h787: data_out = 8'b00111100; // 7   ****
			11'h788: data_out = 8'b00011000; // 8    **
			11'h789: data_out = 8'b00111100; // 9   ****
			11'h78a: data_out = 8'b01100110; // a  **  **
			11'h78b: data_out = 8'b11000011; // b **    **
			11'h78c: data_out = 8'b00000000; // c
			11'h78d: data_out = 8'b00000000; // d
			11'h78e: data_out = 8'b00000000; // e
			11'h78f: data_out = 8'b00000000; // f
			// code x79
			11'h790: data_out = 8'b00000000; // 0
			11'h791: data_out = 8'b00000000; // 1
			11'h792: data_out = 8'b00000000; // 2
			11'h793: data_out = 8'b00000000; // 3
			11'h794: data_out = 8'b00000000; // 4
			11'h795: data_out = 8'b11000110; // 5 **   **
			11'h796: data_out = 8'b11000110; // 6 **   **
			11'h797: data_out = 8'b11000110; // 7 **   **
			11'h798: data_out = 8'b11000110; // 8 **   **
			11'h799: data_out = 8'b11000110; // 9 **   **
			11'h79a: data_out = 8'b11000110; // a **   **
			11'h79b: data_out = 8'b01111110; // b  ******
			11'h79c: data_out = 8'b00000110; // c      **
			11'h79d: data_out = 8'b00001100; // d     **
			11'h79e: data_out = 8'b11111000; // e *****
			11'h79f: data_out = 8'b00000000; // f
			// code x7a
			11'h7a0: data_out = 8'b00000000; // 0
			11'h7a1: data_out = 8'b00000000; // 1
			11'h7a2: data_out = 8'b00000000; // 2
			11'h7a3: data_out = 8'b00000000; // 3
			11'h7a4: data_out = 8'b00000000; // 4
			11'h7a5: data_out = 8'b11111110; // 5 *******
			11'h7a6: data_out = 8'b11001100; // 6 **  **
			11'h7a7: data_out = 8'b00011000; // 7    **
			11'h7a8: data_out = 8'b00110000; // 8   **
			11'h7a9: data_out = 8'b01100000; // 9  **
			11'h7aa: data_out = 8'b11000110; // a **   **
			11'h7ab: data_out = 8'b11111110; // b *******
			11'h7ac: data_out = 8'b00000000; // c
			11'h7ad: data_out = 8'b00000000; // d
			11'h7ae: data_out = 8'b00000000; // e
			11'h7af: data_out = 8'b00000000; // f
			// code x7b
			11'h7b0: data_out = 8'b00000000; // 0
			11'h7b1: data_out = 8'b00000000; // 1
			11'h7b2: data_out = 8'b00001110; // 2     ***
			11'h7b3: data_out = 8'b00011000; // 3    **
			11'h7b4: data_out = 8'b00011000; // 4    **
			11'h7b5: data_out = 8'b00011000; // 5    **
			11'h7b6: data_out = 8'b01110000; // 6  ***
			11'h7b7: data_out = 8'b00011000; // 7    **
			11'h7b8: data_out = 8'b00011000; // 8    **
			11'h7b9: data_out = 8'b00011000; // 9    **
			11'h7ba: data_out = 8'b00011000; // a    **
			11'h7bb: data_out = 8'b00001110; // b     ***
			11'h7bc: data_out = 8'b00000000; // c
			11'h7bd: data_out = 8'b00000000; // d
			11'h7be: data_out = 8'b00000000; // e
			11'h7bf: data_out = 8'b00000000; // f
			// code x7c
			11'h7c0: data_out = 8'b00000000; // 0
			11'h7c1: data_out = 8'b00000000; // 1
			11'h7c2: data_out = 8'b00011000; // 2    **
			11'h7c3: data_out = 8'b00011000; // 3    **
			11'h7c4: data_out = 8'b00011000; // 4    **
			11'h7c5: data_out = 8'b00011000; // 5    **
			11'h7c6: data_out = 8'b00000000; // 6
			11'h7c7: data_out = 8'b00011000; // 7    **
			11'h7c8: data_out = 8'b00011000; // 8    **
			11'h7c9: data_out = 8'b00011000; // 9    **
			11'h7ca: data_out = 8'b00011000; // a    **
			11'h7cb: data_out = 8'b00011000; // b    **
			11'h7cc: data_out = 8'b00000000; // c
			11'h7cd: data_out = 8'b00000000; // d
			11'h7ce: data_out = 8'b00000000; // e
			11'h7cf: data_out = 8'b00000000; // f
			// code x7d
			11'h7d0: data_out = 8'b00000000; // 0
			11'h7d1: data_out = 8'b00000000; // 1
			11'h7d2: data_out = 8'b01110000; // 2  ***
			11'h7d3: data_out = 8'b00011000; // 3    **
			11'h7d4: data_out = 8'b00011000; // 4    **
			11'h7d5: data_out = 8'b00011000; // 5    **
			11'h7d6: data_out = 8'b00001110; // 6     ***
			11'h7d7: data_out = 8'b00011000; // 7    **
			11'h7d8: data_out = 8'b00011000; // 8    **
			11'h7d9: data_out = 8'b00011000; // 9    **
			11'h7da: data_out = 8'b00011000; // a    **
			11'h7db: data_out = 8'b01110000; // b  ***
			11'h7dc: data_out = 8'b00000000; // c
			11'h7dd: data_out = 8'b00000000; // d
			11'h7de: data_out = 8'b00000000; // e
			11'h7df: data_out = 8'b00000000; // f
			// code x7e
			11'h7e0: data_out = 8'b00000000; // 0
			11'h7e1: data_out = 8'b00000000; // 1
			11'h7e2: data_out = 8'b01110110; // 2  *** **
			11'h7e3: data_out = 8'b11011100; // 3 ** ***
			11'h7e4: data_out = 8'b00000000; // 4
			11'h7e5: data_out = 8'b00000000; // 5
			11'h7e6: data_out = 8'b00000000; // 6
			11'h7e7: data_out = 8'b00000000; // 7
			11'h7e8: data_out = 8'b00000000; // 8
			11'h7e9: data_out = 8'b00000000; // 9
			11'h7ea: data_out = 8'b00000000; // a
			11'h7eb: data_out = 8'b00000000; // b
			11'h7ec: data_out = 8'b00000000; // c
			11'h7ed: data_out = 8'b00000000; // d
			11'h7ee: data_out = 8'b00000000; // e
			11'h7ef: data_out = 8'b00000000; // f
			// code x7f
			11'h7f0: data_out = 8'b00000000; // 0
			11'h7f1: data_out = 8'b00000000; // 1
			11'h7f2: data_out = 8'b00000000; // 2
			11'h7f3: data_out = 8'b00000000; // 3
			11'h7f4: data_out = 8'b00010000; // 4    *
			11'h7f5: data_out = 8'b00111000; // 5   ***
			11'h7f6: data_out = 8'b01101100; // 6  ** **
			11'h7f7: data_out = 8'b11000110; // 7 **   **
			11'h7f8: data_out = 8'b11000110; // 8 **   **
			11'h7f9: data_out = 8'b11000110; // 9 **   **
			11'h7fa: data_out = 8'b11111110; // a *******
			11'h7fb: data_out = 8'b00000000; // b
			11'h7fc: data_out = 8'b00000000; // c
			11'h7fd: data_out = 8'b00000000; // d
			11'h7fe: data_out = 8'b00000000; // e
			11'h7ff: data_out = 8'b00000000; // f
			default: data_out = 8'b00000000;
		endcase
	end
endmodule